PK
      RZ�9��n  �n     cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_0":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_1":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_2":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_3":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_4":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_5":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_6":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_7":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_8":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_9":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_10":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_11":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_12":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_13":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_14":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_15":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_16":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_17":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_18":["pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_1"],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_19":["pin-type-component_066283b3-5862-4847-8565-3f3a3ce6a34b_0"],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_20":["pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_1"],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_21":["pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_2"],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_22":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_23":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_24":["pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_3"],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_25":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_26":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_27":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_28":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_29":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_30":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_31":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_32":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_33":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_34":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_35":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_36":[],"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_37":[],"pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_0":["pin-type-component_066283b3-5862-4847-8565-3f3a3ce6a34b_0"],"pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_1":["pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_18"],"pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_2":["pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_21"],"pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_3":["pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_24"],"pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_0":["pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_1"],"pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_1":["pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_20"],"pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_0":["pin-type-component_066283b3-5862-4847-8565-3f3a3ce6a34b_0"],"pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_1":["pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_0"],"pin-type-component_066283b3-5862-4847-8565-3f3a3ce6a34b_0":["pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_19","pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_0","pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_0"]},"pin_to_color":{"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_0":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_1":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_2":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_3":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_4":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_5":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_6":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_7":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_8":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_9":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_10":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_11":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_12":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_13":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_14":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_15":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_16":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_17":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_18":"#ff0000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_19":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_20":"#0000ff","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_21":"#00ff00","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_22":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_23":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_24":"#787878","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_25":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_26":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_27":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_28":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_29":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_30":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_31":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_32":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_33":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_34":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_35":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_36":"#000000","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_37":"#000000","pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_0":"#000000","pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_1":"#ff0000","pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_2":"#00ff00","pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_3":"#787878","pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_0":"#0000ff","pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_1":"#0000ff","pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_0":"#000000","pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_1":"#0000ff","pin-type-component_066283b3-5862-4847-8565-3f3a3ce6a34b_0":"#000000"},"pin_to_state":{"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_0":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_1":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_2":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_3":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_4":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_5":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_6":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_7":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_8":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_9":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_10":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_11":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_12":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_13":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_14":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_15":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_16":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_17":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_18":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_19":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_20":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_21":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_22":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_23":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_24":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_25":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_26":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_27":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_28":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_29":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_30":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_31":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_32":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_33":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_34":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_35":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_36":"neutral","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_37":"neutral","pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_0":"neutral","pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_1":"neutral","pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_2":"neutral","pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_3":"neutral","pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_0":"neutral","pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_1":"neutral","pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_0":"neutral","pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_1":"neutral","pin-type-component_066283b3-5862-4847-8565-3f3a3ce6a34b_0":"neutral"},"next_color_idx":9,"wires_placed_in_order":[["pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_0","pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_1"],["pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_1","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_20"],["pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_0","pin-type-component_066283b3-5862-4847-8565-3f3a3ce6a34b_0"],["pin-type-component_066283b3-5862-4847-8565-3f3a3ce6a34b_0","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_19"],["pin-type-component_066283b3-5862-4847-8565-3f3a3ce6a34b_0","pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_0"],["pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_1","pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_0"],["pin-type-component_066283b3-5862-4847-8565-3f3a3ce6a34b_0","pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_0"],["pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_20","pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_1"],["pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_18","pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_1"],["pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_0","pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_1"],["pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_21","pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_2"],["pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_24","pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_3"]],"wires_removed_and_placed_in_order":[[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_0","pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_1"]]],[[],[["pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_1","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_20"]]],[[],[["pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_0","pin-type-component_066283b3-5862-4847-8565-3f3a3ce6a34b_0"]]],[[],[["pin-type-component_066283b3-5862-4847-8565-3f3a3ce6a34b_0","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_19"]]],[[],[["pin-type-component_066283b3-5862-4847-8565-3f3a3ce6a34b_0","pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_0"]]],[[["pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_1","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_20"]],[]],[[["pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_1","pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_0"]],[]],[[["pin-type-component_066283b3-5862-4847-8565-3f3a3ce6a34b_0","pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_0"]],[]],[[],[["pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_1","pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_0"]]],[[],[["pin-type-component_066283b3-5862-4847-8565-3f3a3ce6a34b_0","pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_0"]]],[[],[["pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_20","pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_1"]]],[[],[["pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_18","pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_1"]]],[[["pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_0","pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_1"]],[]],[[],[["pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_0","pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_1"]]],[[],[["pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_21","pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_2"]]],[[],[["pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_24","pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_3"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_0":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_1":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_2":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_3":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_4":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_5":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_6":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_7":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_8":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_9":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_10":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_11":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_12":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_13":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_14":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_15":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_16":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_17":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_18":"0000000000000003","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_19":"0000000000000002","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_20":"0000000000000001","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_21":"0000000000000004","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_22":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_23":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_24":"0000000000000005","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_25":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_26":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_27":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_28":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_29":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_30":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_31":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_32":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_33":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_34":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_35":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_36":"_","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_37":"_","pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_0":"0000000000000002","pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_1":"0000000000000003","pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_2":"0000000000000004","pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_3":"0000000000000005","pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_0":"0000000000000000","pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_1":"0000000000000001","pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_0":"0000000000000002","pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_1":"0000000000000000","pin-type-component_066283b3-5862-4847-8565-3f3a3ce6a34b_0":"0000000000000002"},"component_id_to_pins":{"c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30","31","32","33","34","35","36","37"],"858a7e7d-4a33-418b-973b-f010608cc0cc":["0","1","2","3"],"399f45d5-3880-4d5d-a7b3-79920b289e3a":["0","1"],"44aa55f4-8b65-4c7b-bb33-cc7d27d3abad":["0","1"],"066283b3-5862-4847-8565-3f3a3ce6a34b":["0"]},"uid_to_net":{"_":[],"0000000000000002":["pin-type-component_066283b3-5862-4847-8565-3f3a3ce6a34b_0","pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_0","pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_19","pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_0"],"0000000000000001":["pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_20","pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_1"],"0000000000000003":["pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_18","pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_1"],"0000000000000000":["pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_0","pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_1"],"0000000000000004":["pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_21","pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_2"],"0000000000000005":["pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_24","pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_3"]},"uid_to_text_label":{"0000000000000002":"Net 2","0000000000000001":"Net 1","0000000000000003":"Net 3","0000000000000000":"Net 0","0000000000000004":"Net 4","0000000000000005":"Net 5"},"all_breadboard_info_list":["bbae4fac-23b2-4c26-9347-1b24e05a4497_30_2_True_985.0000000000006_339.9999999999999_up"],"breadboard_info_list":[],"componentsData":[{"compProperties":{},"position":[758.3564995000004,306.8364994999996],"typeId":"51de4dd0-800a-4032-a9d9-828513b5fd23","componentVersion":8,"instanceId":"c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1","orientation":"down","circleData":[[857.5,485],[856.9180000000001,464.02399999999983],[856.9180000000001,445.96250000000003],[855.7525,424.4059999999999],[854.587,405.1790000000001],[856.3344999999999,385.95199999999994],[856.3344999999999,365.56100000000004],[856.3344999999999,346.33399999999995],[855.7525,327.6889999999995],[855.7525,306.71449999999936],[855.7525,287.4874999999994],[855.7525,267.6784999999993],[855.1689999999999,249.6169999999995],[857.5,230.97349999999938],[855.1689999999999,209.9974999999996],[855.1689999999999,185.95999999999924],[856.3344999999999,168.63199999999932],[856.3344999999999,149.98699999999934],[855.1689999999999,130.75999999999948],[658.2415000000007,484.41650000000004],[659.989000000001,464.02399999999983],[657.076000000001,445.96250000000003],[659.989000000001,423.82249999999993],[659.989000000001,405.1790000000001],[659.4055000000009,385.95199999999994],[659.989000000001,366.725],[659.989000000001,347.49799999999993],[659.989000000001,325.94149999999956],[659.4055000000009,307.2979999999993],[659.4055000000009,286.32199999999943],[657.076000000001,268.84399999999937],[658.823500000001,247.86949999999945],[661.736500000001,227.47699999999963],[658.823500000001,208.2499999999992],[658.823500000001,187.85749999999928],[661.736500000001,169.79599999999954],[658.823500000001,148.2394999999994],[658.2415000000007,130.75999999999948]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[770.3005,767.3735],"typeId":"a983a292-04ed-464a-8e70-77365ceef41b","componentVersion":1,"instanceId":"858a7e7d-4a33-418b-973b-f010608cc0cc","orientation":"left","circleData":[[677.5,785],[677.5,771.2510000000001],[677.5,754.448],[677.5,742.226]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"200","displayFormat":"input","showOnComp":true,"isVisibleToUser":true},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.25%","value":"0.25%"},{"label":"0.1%","value":"0.1%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false,"isVisibleToUser":true},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"string","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false,"isVisibleToUser":true}},"position":[490,590],"typeId":"72c75556-baa3-04e7-55a5-e13f447c8c5a","componentVersion":1,"instanceId":"44aa55f4-8b65-4c7b-bb33-cc7d27d3abad","orientation":"up","circleData":[[452.5,590],[527.4999999999995,590]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"HLMP-AB75-WXBDD","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"Broadcom","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[549.16975,508.29275000000007],"typeId":"88687a1b-2b49-a94f-aa87-8f037dbbcbbc","componentVersion":1,"instanceId":"399f45d5-3880-4d5d-a7b3-79920b289e3a","orientation":"up","circleData":[[542.5,590],[557.5045,590]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[317.350642,693.43517],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"066283b3-5862-4847-8565-3f3a3ce6a34b","orientation":"up","circleData":[[317.5,665]],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"109.17577","left":"282.19617","width":"648.10433","height":"818.19773","x":"282.19617","y":"109.17577"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_066283b3-5862-4847-8565-3f3a3ce6a34b_0\",\"endPinId\":\"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_19\",\"rawStartPinId\":\"pin-type-component_066283b3-5862-4847-8565-3f3a3ce6a34b_0\",\"rawEndPinId\":\"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_19\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"317.5000000000_665.0000000000\\\",\\\"317.5000000000_484.4165000000\\\",\\\"658.2415000000_484.4165000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_066283b3-5862-4847-8565-3f3a3ce6a34b_0\",\"endPinId\":\"pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_0\",\"rawStartPinId\":\"pin-type-component_066283b3-5862-4847-8565-3f3a3ce6a34b_0\",\"rawEndPinId\":\"pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"317.5000000000_665.0000000000\\\",\\\"317.5000000000_620.0000000000\\\",\\\"392.5000000000_620.0000000000\\\",\\\"392.5000000000_785.0000000000\\\",\\\"677.5000000000_785.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_066283b3-5862-4847-8565-3f3a3ce6a34b_0\",\"endPinId\":\"pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_0\",\"rawStartPinId\":\"pin-type-component_066283b3-5862-4847-8565-3f3a3ce6a34b_0\",\"rawEndPinId\":\"pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"317.5000000000_665.0000000000\\\",\\\"317.5000000000_590.0000000000\\\",\\\"452.5000000000_590.0000000000\\\"]}\"}","{\"color\":\"#0000ff\",\"startPinId\":\"pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_1\",\"endPinId\":\"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_20\",\"rawStartPinId\":\"pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_1\",\"rawEndPinId\":\"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_20\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"557.5045000000_590.0000000000\\\",\\\"625.0000000000_590.0000000000\\\",\\\"625.0000000000_464.0240000000\\\",\\\"659.9890000000_464.0240000000\\\"]}\"}","{\"color\":\"#ff0000\",\"startPinId\":\"pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_1\",\"endPinId\":\"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_18\",\"rawStartPinId\":\"pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_1\",\"rawEndPinId\":\"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_18\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"677.5000000000_771.2510000000\\\",\\\"640.0000000000_771.2510000000\\\",\\\"640.0000000000_545.0000000000\\\",\\\"887.5000000000_545.0000000000\\\",\\\"887.5000000000_130.7600000000\\\",\\\"855.1690000000_130.7600000000\\\"]}\"}","{\"color\":\"#0000ff\",\"startPinId\":\"pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_0\",\"endPinId\":\"pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_1\",\"rawStartPinId\":\"pin-type-component_399f45d5-3880-4d5d-a7b3-79920b289e3a_0\",\"rawEndPinId\":\"pin-type-component_44aa55f4-8b65-4c7b-bb33-cc7d27d3abad_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"542.5000000000_590.0000000000\\\",\\\"527.5000000000_590.0000000000\\\"]}\"}","{\"color\":\"#00ff00\",\"startPinId\":\"pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_2\",\"endPinId\":\"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_21\",\"rawStartPinId\":\"pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_2\",\"rawEndPinId\":\"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_21\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"677.5000000000_754.4480000000\\\",\\\"602.5000000000_754.4480000000\\\",\\\"602.5000000000_445.9625000000\\\",\\\"657.0760000000_445.9625000000\\\"]}\"}","{\"color\":\"#787878\",\"startPinId\":\"pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_3\",\"endPinId\":\"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_24\",\"rawStartPinId\":\"pin-type-component_858a7e7d-4a33-418b-973b-f010608cc0cc_3\",\"rawEndPinId\":\"pin-type-component_c18bbeac-df6f-4ddc-bcba-5fd80b7ea1a1_24\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"677.5000000000_742.2260000000\\\",\\\"587.5000000000_742.2260000000\\\",\\\"587.5000000000_385.9520000000\\\",\\\"659.4055000000_385.9520000000\\\"]}\"}"],"projectDescription":""}PK
      RZ               jsons/PK
      RZ��       jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"ESP32-WROOM-32UE","category":["User Defined"],"id":"51de4dd0-800a-4032-a9d9-828513b5fd23","componentVersion":8,"userDefined":true,"subtypeDescription":"","subtypePic":"61f598ae-58c3-4b7b-a0c5-99e4be3565c0.png","iconPic":"b240e25a-70ca-477b-8a45-be7a3295a83b.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"14.24371","numDisplayRows":"25.02143","pins":[{"uniquePinIdString":"0","positionMil":"51.22883,2438.82817","isAnchorPin":true,"label":"3v3"},{"uniquePinIdString":"1","positionMil":"55.10883,2298.98817","isAnchorPin":false,"label":"EN"},{"uniquePinIdString":"2","positionMil":"55.10883,2178.57817","isAnchorPin":false,"label":"VP"},{"uniquePinIdString":"3","positionMil":"62.87883,2034.86817","isAnchorPin":false,"label":"VN"},{"uniquePinIdString":"4","positionMil":"70.64883,1906.68817","isAnchorPin":false,"label":"34"},{"uniquePinIdString":"5","positionMil":"58.99883,1778.50817","isAnchorPin":false,"label":"35"},{"uniquePinIdString":"6","positionMil":"58.99883,1642.56817","isAnchorPin":false,"label":"32"},{"uniquePinIdString":"7","positionMil":"58.99883,1514.38817","isAnchorPin":false,"label":"33"},{"uniquePinIdString":"8","positionMil":"62.87883,1390.08817","isAnchorPin":false,"label":"25"},{"uniquePinIdString":"9","positionMil":"62.87883,1250.25817","isAnchorPin":false,"label":"26"},{"uniquePinIdString":"10","positionMil":"62.87883,1122.07817","isAnchorPin":false,"label":"27"},{"uniquePinIdString":"11","positionMil":"62.87883,990.01817","isAnchorPin":false,"label":"14"},{"uniquePinIdString":"12","positionMil":"66.76883,869.60817","isAnchorPin":false,"label":"12"},{"uniquePinIdString":"13","positionMil":"51.22883,745.31817","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"14","positionMil":"66.76883,605.47817","isAnchorPin":false,"label":"13"},{"uniquePinIdString":"15","positionMil":"66.76883,445.22817","isAnchorPin":false,"label":"D2"},{"uniquePinIdString":"16","positionMil":"58.99883,329.70817","isAnchorPin":false,"label":"D3"},{"uniquePinIdString":"17","positionMil":"58.99883,205.40817","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"18","positionMil":"66.76883,77.22817","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"19","positionMil":"1379.61883,2434.93817","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"20","positionMil":"1367.96883,2298.98817","isAnchorPin":false,"label":"23"},{"uniquePinIdString":"21","positionMil":"1387.38883,2178.57817","isAnchorPin":false,"label":"22"},{"uniquePinIdString":"22","positionMil":"1367.96883,2030.97817","isAnchorPin":false,"label":"TX"},{"uniquePinIdString":"23","positionMil":"1367.96883,1906.68817","isAnchorPin":false,"label":"RX"},{"uniquePinIdString":"24","positionMil":"1371.85883,1778.50817","isAnchorPin":false,"label":"21"},{"uniquePinIdString":"25","positionMil":"1367.96883,1650.32817","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"26","positionMil":"1367.96883,1522.14817","isAnchorPin":false,"label":"19"},{"uniquePinIdString":"27","positionMil":"1367.96883,1378.43817","isAnchorPin":false,"label":"18"},{"uniquePinIdString":"28","positionMil":"1371.85883,1254.14817","isAnchorPin":false,"label":"5"},{"uniquePinIdString":"29","positionMil":"1371.85883,1114.30817","isAnchorPin":false,"label":"17"},{"uniquePinIdString":"30","positionMil":"1387.38883,997.78817","isAnchorPin":false,"label":"16"},{"uniquePinIdString":"31","positionMil":"1375.73883,857.95817","isAnchorPin":false,"label":"4"},{"uniquePinIdString":"32","positionMil":"1356.31883,722.00817","isAnchorPin":false,"label":"0"},{"uniquePinIdString":"33","positionMil":"1375.73883,593.82817","isAnchorPin":false,"label":"2"},{"uniquePinIdString":"34","positionMil":"1375.73883,457.87817","isAnchorPin":false,"label":"15"},{"uniquePinIdString":"35","positionMil":"1356.31883,337.46817","isAnchorPin":false,"label":"D1"},{"uniquePinIdString":"36","positionMil":"1375.73883,193.75817","isAnchorPin":false,"label":"D0"},{"uniquePinIdString":"37","positionMil":"1379.61883,77.22817","isAnchorPin":false,"label":"CKL"}],"pinType":"wired"},"properties":[]},{"subtypeName":"OLED 1.3\"","category":["User Defined"],"id":"a983a292-04ed-464a-8e70-77365ceef41b","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"9bab9bed-0662-4eeb-a3ad-16a556afeca0.png","iconPic":"0291db46-fb1c-4fc7-8f6c-e1e807286f19.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"20.00000","numDisplayRows":"20.00000","pins":[{"uniquePinIdString":"0","positionMil":"882.49000,1618.67000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"974.15000,1618.67000","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"2","positionMil":"1086.17000,1618.67000","isAnchorPin":false,"label":"SCL"},{"uniquePinIdString":"3","positionMil":"1167.65000,1618.67000","isAnchorPin":false,"label":"SDA"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Resistor","category":["Basic"],"id":"72c75556-baa3-04e7-55a5-e13f447c8c5a","subtypeDescription":"","subtypePic":"bbfae99c-8036-4c5e-89fd-a87441410720.png","userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[{"type":"double","name":"Resistance","value":200,"unit":"Ω","showOnComp":true,"required":true,"validRange":[0,70000]},{"type":"dropdown","name":"Tolerance","value":"5%","options":["0.25%","0.1%","0.5%","1%","2%","5%","10%"],"showOnComp":false,"required":true},{"type":"dropdown","name":"Number Of Bands","value":5,"options":[4,5,6],"showOnComp":false,"required":true}],"iconPic":"a262aa33-74c4-460b-b0ad-c746896f6744.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"LED: Two Pin (blue)","subtypeDescription":"","id":"88687a1b-2b49-a94f-aa87-8f037dbbcbbc","category":["Output"],"userDefined":false,"subtypePic":"d8ab57a1-5a79-4c55-bee7-02b60939cb6a.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"62.87000,0.00000","endPositionMil":"62.87000,-341.89000","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"162.90000,0.00000","endPositionMil":"162.90000,-341.89000","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"2.14670","numDisplayRows":"4.05650","pinType":"movable"},"properties":[{"type":"string","name":"mpn","value":"HLMP-AB75-WXBDD","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Broadcom","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"cc0ca695-66e1-46bc-a2f3-28706ce884b5.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]}]}PK
      RZ               images/PK
      RZuA�V� V� /   images/61f598ae-58c3-4b7b-a0c5-99e4be3565c0.png�PNG

   IHDR  ,     F�t'   	pHYs  �  ��+  ��IDATx�<}	�\U�����[{�����tV��$,*.0��#����8�8ʀ3#���<n���  ".��!$$dOw�Nw����ګ�~��~��ԃm��ܳ|�[�o9����%U!��@��e��}�E1
� ���(��o%]sG�e��JU���˲2�&۶}����Sooo��:�7<�X,����Q�44F�����"A
��n7*�Z�TJ�$I�X~��)�'�=HN��4zȘ�\�ā��Z�R�V㉘i��Z}FA���	���(���]����a���i����^���&�$�=���
^�l�A��&��\��躵ZMQU|�p\L�0�hY��0C�����ҢH�����h�DU�D"�Jԉ��X:�S�g��s����sUS���	=�ȦQ�����t:����`\����5]�C�f�A�x<�x��э���<��h��2���H�������Vв�k%�ej~|ff&�Ȃz�RÊ4Mǎzϴ�u`n�Ek1b*�z&�Hf�š%��|,��̆oeU�襠}L3@�r�����D?�\��b�������U�g�0"ʈ�����s�cM���-���U='���[KThΉN�Wt�LU�_Y�v%��8�^$I��:��m��	�"+���a@lۥ��$?�WR(�*�j��$��<Y���@�l��U�W44��4u��Wu��H=�� /����~��}���%)�ȸ�$��Xh��>6�X�vvv��?y����ß455����l.���陙�(B+���;��*�x��܌ަ�
 �()`��(��˦��ƈ��*�kv\��/;u��hym�_/
�ځG��l6��;w��Mc�\�n�����"�X��T*%�!���d 7��TD'.	Ct�q��d �iɘ�.k�N!"��d	Oɒ�������6��-h3PFW�������}/�����Y�s�?���R��1kb�$r>�����O�q�b�T�lI�$3tmbq��E�*1!�?�[ݪ��1[|�o��|��rY�$�#x�E{�&���['�˭��׭���	Iijmm]��b�t�u�e2N3"=뺉�A|
!�/CR�k���A���$h
�EY³��*��BHS�,��$�u�BR�`ZUum��Dڑ��|�XDK�>xc�$1f�1����vp΁z���y�	�,zH�q�"��&+D��N�@O�OA����+����lAWG7�g�i���ޙ�d
�2�%�}]&��i�U#p0þޕ0�Yn�eW��d�(����`�C�B"�3�<��?��/���L
�@��B.������Ek�LOO��֯;r��X1]K�V�H��ݽbŊU��A_6�K]�=M���'�Y�eSiA�i��ibe���mmm5���`���%�kߵ��7�������P5BX?)>�QbB0�W����~������W+Woڴ	\� qMMA#�Huih������]BX�z��m$�N�t�2�`�/��$�0~rbF�*���$�\U����~$`�D����ȅ��%�I���܂�!�3*Sh�G�'����)
Yl?����W�`Z�Nʛl��s��ْ���B�o��d�i��O04!�L�?�We�0V��FN�=����X�b0a�N��Z����(��SD(.�$3�I�CHJA�i��ԃփ���Ob��$�CN�����H�d��,��C����SG{]�@4�#Q@�o�� $���$a�#,V�-[�ޭ7,[�����/��;V����L��3�M�X����<�) g����L��,��V#��T*y��qҧ��P�`~�U�q�X,3�'�H	HE�)�d��U[�l��W�D3TXw�(G���%3i4�����?��^�����+����qSE)���!1}��������>��O��k�o	�\t뭷>���`#7m^w���
�4?;��ח\�bdd�C0`��5Ab1���w��n�_�O|>6}
�;���l�I����W_�|�ٳg�u�4���s��^z)�.]�P�u�E�ʹA�z�XPf���9��$�F��Jl� �]��9<Ga/R�
�C�����!�H
B��.$�n�X����1!8��X
�[̋��&@�"��#���߆� ��&�``��BK0�d��p�h��"`ϒ����˲�o�L`��$୩�p �|S4U .�߻�����^�Z<�CŪ�=2������� b��v�B�l�X���TBn6�/WI�
\�O���T�Кe1P�δZ�A*íq�B��'��W|��T��q�@��r6�RII�>����ɝ���D�>|�.���ʂ������tX2H��W�\�����A0g<^��@��}"�����@=��ϢMi��A�LU��_܉���˟o������C0��%(@��\�����܆=�x�4� ���l%S;�Ǆ`��{ڎ�:;;;}�Ё͛7^}�Uo��F_/�玞9��+o��=��w�q���i؟��6�߿�R����ϼ��k~��~�k_��c&�W�O`�����%�S�d��$K�
��3��#W�Q�ZTY�Q�I��������� E�cǎ���=�<��������X: �,����D��8��\;�4�퓩"^� ���	M
=����N��"K��&�%ؘ��+���<�@����0�����Ln	b���e�P+<P�eq�
���$�J\_>/��u�+?j�	�g0$��-z�fj��\(.�D�M��3ς;�|IT���Vڜ��ɽ�I���C������^0�8ױdAc�G		@�@�i���(@�a�C��C�X�&� �实eXR��0��p�ّ1� b�9��&k�����T�@�8\2hUX��
��2,NM�$rS�K��8�>Wk����DZRO�.���vŮ�rx
k$�I �7t�W@��M�OC,oz�?B�7�ӗ]�uvf��_����U�O�Y�jd������t:�G�^�@�ح�۷���}���x�7�������C��~�C�����v��E���T�~������[�n��A�@g�^�
=b�A,X-=�!Ɋ5��O��#��7�p�#�<��&�<`ϣ� �3�����7�ӟ��?�V`� qx#�4���ò�o��S)0zsg?Ĳ#�b��v�� �oq7$����aWո���{���?����~�{ߋ�F�+�0C�0�
�۱lf�� sۥ).¢�ŵ$Y�����Nœ��� |��Lx�C&2>����0A;�%xdbj��D���W�y|+I虋%zf�����A��"��ӎD����ur���· uÀt$���VmԹ9�2�m#�` �CC�7�,Gڽ^���09��՗�oo���n��H�<���qb�
�Z��Kꀍ��_E�^dm"� 	�`�1\*���,kX��Fo 2vAS�h�;��sG�B_,��u���J<�[�N��
]��x=`���/~񋓓��!���Z���Uk�#G^m7��L�m~��+���W���B�H�R��|�}7�w���_�ϻ�!�!½�X�D#� Ϯ\
,(x>��|����{�|���G?Ĝ���o�k 	,�J�ȇ�,�$�.����A�TXp�Z9��[�hQ"?x�`�L��okn�<��sss�u���n/m�S�t��xP\����Pߢ�T6WP��C Z��O����������}�z�ٌ��#�$�S'%/[�.(Q���	��|�� �-��G��+�V�Z�f͚S�C�D��W�V)��U��"%�-�p��P���n��Ʉ��n�V�XⲄ7h& /4cxOp=/?7�b!W�o��f�w�009D,�*+��R%Q:����)��G X|E�|�`�y�H�r[��?���ި�7L��lΑI����#�Vd/�Hq4trө��g5nI#���5U��x������5Mmm�x۵z�}鍋.Z�I%ɳH��y &����H���{����0�4�fS<۩۵3#C�m�(2��%�؃�%IU����cղf�i!�[��#�\VP���R�x���׷��|!3~��r�*�p���ۼ����B�Oa%L$���%������ݳg����s�ή�|�{�%�������������ޯ~�K�Ї�y��{�ɦs@��I�(pnrbɒ%����׽�:@q�h�<�d���"@�Wv�t=���?��O�������Kss��M
�����߻���>��Ç���.��z���-}F��'wvaa��Ű�h���O�81To����\�N����������w^W�{��n���Bs.��Uձ��n�
������{��ގ�� F���&�`���	h�y�X�.s�o����z�����ꆲ��<�h���gd�B��i�L�,��<4�M�$�C�����{\�xh��]n�8˂<���[rCG)���ٱI����J
8,$|*���	Q�ϻg�(q�QS.x|��At>$3�Vg�[(�#���/�'-�7�J\u+���ET� 2�!�@��yL��5�9y�;���s��-^܇��@4�4�+��(.�SDZ���Ne�,z��� ��aY,2F���� �`�x*��#� ��l� K`k'�x!�D�z���V�l,3�2������q��1�x��f�>����y̧2U!>d�������+!c@y�yfz�37�k��8�Of2��t���[�¸��ioo��Y���A��u�]w�%�8�X��-�/�mc��-[d%��d��
�� &V
���������}�|K[�/��;v#eҹLVN%� Y~v���[���\l������?�V�M%����K:���~宻�^	p��o�0�۷_
�ٵ��������N�u��P�����?�����o~��x*U�ֱ)`C(��D\��[�	����߈A��������bsj����s�������B/����f4Z�K&�rkB�V�^H.f�yR�Bn��P-�6J������g�T� �JPG#SGh�Ƈ%�� ��ÿ�zJ�F�,1L��0"�9	������x��ⱺ�Թ)�$��)`��1o��Qul� �>��b���I)0s�pJ1� �sf�5��ɦ9 �����L����V/{%/�J(1��|�_���?�����P����m{^��ѣk׮Ă�2,�^�G��u`�p: ��U�U%���n #P�	v�Q��=[7�(�|�Ig�~`���]�z�B����!GWL Q��F�}^`yE��b�*�����׳v�Z-�������B �Yv ԑ��趽����\�B�RZ�����寊E0$@b�R��	Q����Wk}��*���X��\�f������� ;�jP8���򮮎ض믿����鑑�l.h	���Ĉ��r��_|�5�,^BA�6��)0��W���|~z%����K,Jj9r��J/�$�1�
]A��[B�}��0������?�;lզ�A�|�9�j�#%=� P�M�b�Q⸍�}Q���)� H`������[��?�ơ��9��صT��X�f�"��� �nb����o�gϞ��'��Eqzz���<555��`o�#��LOnw�䏧�8�+�g|B���`���TȽq�� c�;����X�D"�7��,%j3�FU�
�l����j:�'y(�����l4"����?����i�Y]����r����+�X��Q�!�.�GQw)��,����L��c���\�3����2�N #�ٙ3g�$�=�
�2���7X�j��]}l͝UB�D1�y�i��H�(����%�,�,�>�)�,?��Ap�Q,��K/�vL((���%�Y��2~��{�ԜL��s`E�:��:�S'w�w�I.�� �9z�[����z�a!�ϒ=�1���}o�:u*�L����v���!�@]�~������o~�ܹR__��� T�,�w��\��\�� ��*H[[������m�
J� �X�
�ݪۛ6lx��Q��1���P�_�b��/g�3���z�O=�O=���Ht�5c��2yw�dVS�[s�q؎�p�~�� ���aB�N�ĉO>����ɭ�fa�'C�d�Pҳ�x<�I��"-(ǪQ P�zMǻ0�d�4u�:�e�a��^A격4�P�UA =8'�e�|b��~�d�I �O��X��%�!�<�A�Q��݈���R��,UG��-���P�N�%�=2��`�a(J	�=�3��3�=�i�&	�[̣��X�P	�&M7�iebVE�Lg��R$,�kJ'���e�<Zk�}0���P����Z*�����ī�� ���O$̿��E�]˖/�[�?���\;��=;^��}}���
se&A%S
&yP9��\���e���%��R��^�fx�� Z����TJ�����p8д�3��'l�)����~˦@�%oګ��:2jN�����yG�l��{����W���CaE��J&��Y�i=&_u�eWn��ۢ,�$�z��~�Ԝ]�|���5Sq�g.���%�p^��x�����ܝj��1-���Q�� ��b244	��ܜ��Ғ^}����������A�Y�[��T>E/+|��f���\�(�_�����h���������0]?R�$�/|�c��wC_���w��O>�bŊ�"�uww;.�E��,X��|�3���7'S�8_�o�����뙅�˷oN�.F;|�C���)�na���6��l?&�,yGg��	yb��GP��f��݂͵,�R�h�F�݂i,M|!'NBYg�&�܈11��x�4��9�$��%SI����8��Q>��iIxhܞpKH~�p�!�gꜥX0%��G�d��Tږ�%�̩L��{ 3M�/�a�L:�榨)���H�2i sM�m2٠�8�^8:�:�����j͘Gǳy�G� L�#���+h�Qv��bi�d��7�|�R�t�SEؖ)V����fe��d�Wb�	�$����ru�a�z5���kv�=97Wj�E����僶��q��|t���^�����{r?$�1�'T^&I�x˄����9;�|�J�j��-̬E��3	����!��_�U,T̤(�������'>!�}�����h�D��?�h۶-X|̌	2<� ���LM��a�	��
���^���^{��r���5~��<oXE�E�!��i��x�;޺nݺl�铟��۱��R&�	VXhC�c��>����t*A���)�:��`���&_/��֭�wL���.�I��ˍ��̠Q�xP�R\.W;�H�
��0��)8��J��"�����	߫C�*��3�DEX<��e5�1�IU"�
��O`H*��JAJe�؏��z�y�7�TXuV�7xA0G�L���R�Z(�9n�,)���}*�4,�B)�ɰ:�
��I5�E���K��y}კ�s%хQ&�A�0�N�������.�l�&�2cn^���z�Oa=���Mt�Ōx"%���B�v��nR �a�ڣ��M����\<^��Jf���f�
e��:���H ������fݺ��J#ib/	��qn���okʁ%@�R� x�)~
�P����HE�6)�\�)M�l9H�T*�l��BW����\�K����e����aI�R��`�[�6ƴ������c��z�q�,"Mmי�`���Cs�������/�B86q�X\����G׍]�_ݳw/��Kޒͥ��S�-�&{�Y���1�Q�V�48�ai+@[��g�}v��=�@�U`��Ύ�FC���:0��c�.��y����;���[���_�N�IP~��C��>������:�M�kn��-L nP$
#Fs�1~��'1+��(��`?�3q}�>�e�~r�0:�e�еT��(�4�|��I��L3�fT
��^�>0Ȋ�lܸ���/a�d
��T�R�I(rǆG/�f��R�xP���Bv�Q��{�L�di%�E;�GDt�.����Y�ʛ{ r|����J����*��|�I�U��b_�mr���#��r�����X>_7�����zi��%�R2��}?�2",������������᧞z�Ri`,a�����O>.AA�
t1��H�E��\<�Ol��Ө��=\v¸�}�@y��6��bw�2�/�ϗ�PA��́&矰 AV�y��r����D�09�(�T��U�9�B'z�
yx�j��Ƚ�����#~�>v�ՔBݗ_���=����x����̋������⩫��jfmjѢET\�{���k_����(�S�Y���_��]�^v��s���@Le:?}�Ё�s��S��O?�4>�]X(��b8~v<������UQ�!H�6^���ߪ�������ߎ:
k)��q�e�];_y�f���u6nZ��;&	~:��t�
O*�W�`�l5_
���Dժ�2_L�J 
�Z�SnojN�;����9��
-����z̄�min���Ö���w��'�0]5��Z�!���'Ϟ�!��l���W.[�b�˻�����l�@�CrBBd� ��4�.�mT���B,QUi�
�I�E����*��V�Xf,.�e�9�J=b�&��e��'�XY��2إ0��`#y"��p�-7`�@Ԁ
m @�Ut<�6ay`J�$?�����1mnnV�V��(e�x����,�1���Q$RQ �K�$�0���ް�X�f�/������U��@LX��0��� �~p��,�A�#�l e��"h���Ӱ,�d�X��H�]�{v9nJ���7o�,Ⱦ(�8���F[{;�x||^��E�l)8E��ڙLnvv�|��	|�x�a��Պ�b���B}�ܬ�n�TC0C�� ������q��Bx>���
�c>��81t����3?;	e�lp�L$�>������;!��K���=8гX-�\A�>��3���W�r�UW�ݛϗK�j�)-0��*TuJe�X��h�A�v�fh I^X ƅ�#3e��ޞ01�K�D�,�}�a�%L��ӧ1{r��{���1_ �)]��ࠕ+W���Ǐ�CCT}Wy�D�h�
b P��\rI�Jɍxl�� 6TL�Y(&L�R
�}�����0P2�Q8*Vd��+�[���^ �lش���9Xr�1�993�]��/��!U��p��}� �CR�	�*7z,]qރB�Ʉ	����d�&?R��|�в	V@�p��-��t`*���"�u%ђS�G� ��hj��<�I6M1���*<'A�̘B�/�pl�4�'�H[F�4vʁΎ`��Ep�) |�%��ӴjJ��K�p��J�s�N��@K��M(/,dn~
�c��!�`6��H��ucnl1&�t�2�ĔXL���?�y~ffٲe�=t���9���A8Ewl[����^��`	�R���A�-O�_�Ha�+L��ɓ�ׯ�Tڮf�:;��8` �`$3���[�mf3�a�l3Յ�?��/��)X8O<�����]�o��K蜍D� ����_@t�,��s���0^����6m�����:!�Xvۧn����v������)�ӖJo\����SXX[[K&a�ۻgĩk�\ݶ�;��4N�BĠ8������;�z��mo���)�*��ɉ�Gy�ؑC PϢE�P�0Cۙ��93
�	����<<|�{��A�+-����jQ�Rqx���]}����%g!�%��А5�;y������=����Ix���-���vT-6T8���E!'���b��}6�P����U�z�V�'�K�-�,�eMM�)�,Z��,^�T��G��p)#�~~������=��X�J��f�ĉn�w��-����KE�?dᓗ��^��Ꝕ�c$�<#1g��f���,^�p���8~l����2�,���|��=����wBqa�6��F���~C�ݸ	���K����+���o�.���������nwbh�� ^{�*�'��*>���,[e�̢̦��.zj�y`U��#���OJV芺��M=�LIɡѡl�*r�Q�E���6�sr�X�b��ͭBߒܹs��q�L�Z:p�@�^�bb$)�L��N��P�w7�dgg'�J,�7�Z5"�U�g�m2:<�c�O��9�)CW�a5�̤�d&9T�?��8ۚ	�&9P,�o6�%7�ې4)nf_(T�#HK)t1�t|�����[���)h�W��k�ΝP1k׮��K��b	�ڨC�RX{�J�_�Ǌ$���S&;=#�������o|��Ǟ��$s-� ��_��h�n�����w��!h�K/�������&�/�2���Ç�_�=6����{h,Hv�\eg?��O?������(��⋷lݺUS��رc��]0\���:�e$Jু%�Я�,6:���	�q����f���4`�?�O��?��������*L�N�(�I��8�9��,f�N����9��Dxzk7]>~}�(�W-���k�֫9O�Az�����^�-9:A"�P]s��X5�6�M���cp�"�񅠧�G1C�sUj����Q�r�)�ĲS<�֫5���}�".G��:m�"�!�bt�)ײk�.h������8����<�?8x��q<��*>d�
��L1�ReV��KIA�7hqh�-[���TKiS��rU�c���ڂ� ��vI3`�h@6�|'�X�cM����������L��z��#�T�eϗ0��%�jba��_|�}�	+��"���M��5Պu��`�TE+@���(�JtFԷ�b�;��˲�12��j�{��]{`�s�u�\����射P@E���E�2Ϝ0�h6�~�g�nXF*%���_��3gF$��� ����9t+Y�`�	�]u���Lt{��+l�q�:8�V��"l%����=��c�U����c��Í������P<�T��������<��yh�`��:�=f1��LRz�w���|��w��]K�n��p��s�?�m�\+�2�
�;/��+W.��O~�\�ֳ�l��z�E�'��Ov4M���5����'Z����n��y}��-m���%�Z<�۰��� @9�y��)����kA�p:�ׂ3���X�[L�;̩�B�8"2�xww�a�`�4������<dX�?7^$R���%?�K����=?7BG�)�?r�K{ 6;��L�*��"Q�V)^E�D%�'���R� ���2ȫ�\C��h/��
s��%]�q�=
k֬�b��pb=ǋIb`Si�&FrD�ԡ$ڍj_O:i�&�����V���:9��=.�tܙ��Wʒ�	�N=���V �C�ޜ��$Q�K�,1����I1�����S����̺5+���k��c1��&/���&O��Ĵ7��4�3��D���x��j�������ǰ�d3�g3FU��ԓO>�����vɆPk��RRx�h��5�~�HP��R�!�Nn���|y��CK��ںmn��+m�}[��n��� T�O���5�\#��n�Jcu�6n�pՎ+�����|�_��$b)��/���o{|b���v�+�O�%�P��wQ*��lCe39M~��(ˎ���˦� 9{��1==�Lg�<�3544�mŊ�����`�WTEa�CUh/��3�D�=657�(KLW����+�-��2@�努i�
���Yp�b�+�V���X|��M�`]|����=�>��3���N�vZ��o�LJ̄޽�Ə~�����ӛ�; oK
�y^�T�N��W^y�aq:9���?�J�O:�Ī=B�L!� c�g!�����L:M4yr�4��ƴÐL$�"uR��
.C\A���P�N�7���	f�0"�q"Q�Q2<��!�Kz� �����Nr��]�ۉ��5�
�F0:/\�C���T&)�� 5`w��`D��T��!~,9��A�t6��>1g~aj�@�v#Yg�R Yn��e�(��GxlzlL
�Y> Xd��YZ(P��L�� >��z���e�<��?qQ�m
HS��$��$�U��
t�:��bNB���w�sad@:���P��PYOD��\��Q	��y�Ǟx≬ڄv�[=u��멄mp�i|���w�s�=��w���w��e��������&4"�jX����.ʬ6=A�PT9A�L�Y�y�޽���۰)`~,v�.��_����ݻ�PسgO�P������+6+�4l�$(���_`��u@O�-��X�L���y���PF��kNz�?�#(�������0%�ήU\ˮ�����F2���D�c{p�:{;A�l�7�$�ʡEМ�AWmȠ�n5�t�K�A�Rh���g�<|&O��X��;��W����Qs�{0"a���v���BS3`�iؒ�{����A� GA\
-i��A��B�c�|>���W_��cn�y�����M���p����B)���������/a-�moܸq�Uۉb����vLWF��`PX��.`�F����S�V��egғ�e9=�f�L��=x�O>��v���촩�ڦ��%��c������*
���T��9{� �U^z�]�^��R�ᡣ2�U��	at?H�0
���J��G~u���3#��}��Ȗ"����_8q踪--�'f��s�O�W�_^��X��秧�?L(�k�7���072��(GhD�\n++ڎYu��2�����9��n�����Z��B�D���������/ٳ ���v5�wGO�j��J�-W�y��o�~���{��s��\�}��ߓ�;q�b�3��m����_} �p|�&�lc�e�ﯿ���A�q��=��~��0ǎ��$���|��	��:7���]��3X��K1�;��BxI�.�����B�Ѣ0'�%��%�5e۶m?�����o۶]��o/�z�B�0YLRE�a�@�%����ߏ?��C���-�|Ω�����������w~��?f�M(<.�% c�&[�!]��At�(���-Y��k�C!,^�K�T�94lL"&ּ��Z���'F�����X��)�q��z&`�C�=}��RGgW���ˇO����֎�c8���t�0��W���P<�ơ8%?k�"I���6d�C^p�V(�o�<��	/U�U��A`�h�MTH=�A)��pE��xO�+X�Ut�¤����B��Ux<�I|���$�i^6��f0���4A�FyE�
�b"!p��ň� �����6r�(�&'�xw/z��[g�N�ڶ�uݺu�'�g����A�޶n�a��k�2�X�'y1Z:b	I̐i�`��j��w�y���k7=5&�*0�[VQ'	��5=����D�}�u��c���z�'P؟~7����ӳ������h0 ���G�<���tu@��{ｿ~�G���I�c&o˵ ���G=��݁���`�Z��u�9;�>�sh�v�Jt�y���}�\r�% ��u��
���ỳ|���g���[����I�L�s�v`����¼*���*���j�N)^�D�� ��_���ۿ��w�� <o�� �v�&$����^��AS�t2��L�3�HZ ��9����WX�8|��)R��Ե�c�+֬�TN�N����mikmnk�h5�F�9��|��r2��UV����I<��4�.�c{�
�tWJ~G(P�`�L*Sg��۔�]�˼(���J�]��;��Э�P���2��
ˣq!L��Ǝ*"?�#��j���
A@V�z����4�0m���/�����9��	 ������9|�e@P�<��Ű���`���^X��,:�@���<��CY���C�g���2M5zT��"��YJ�ӕS�t}�9�^ܓE��r���#��i#�T�u������p�D7�9��)x�՘.�^^�"�+;�t:?��?}�T��>���Q
�Z�%�*co50+e��J�5m�9��J�Bvue��+���17P�s��#�{�����'f�A�zCTդ/V�Ƚ�����ڨ��$$��S/�ݝ�	3�\&�ڛ���-7�����7����������-r,|��b#~���SY�q��� �-[��$8���c��oxo�x"�`�\P�b��M7ތy�S	�����)l���e,�)�k�n0�TUEE<(DwťR���z��?�8�$��� H
˧��<1ld��8,��D����w�m߾���݇������mٲ�'�
mzzz�m(pC׽��y������L/�=4��o���W���)_A.h�}.L�۪3yl9?�Gg����oTA"}/8ܔ��Y��<}����-�Ǡb��P�d<ūC�9]����r*8]�6m���H�
�)bY���^X87�5�� �U,�3.{�g��-���lt���
��ȑ#�d�Ӑ'$�o��chf��~�?p�P';=��x:�������4y����1���֠[y@@�+@QX0$�Ю�Ѝr�Ba�EP%�O����"�V�`�r���TY�?�l�2�]�R?��Ӡ@{g�^�>�М$�l�R�С�c�uua,8#����:;��H��&"�HS�D5ON��v�����������{9�@
~�gh��0]�����z��n�y�E�O�>��xVķA a���b�@W�����l�OQ��ߝ��o|���ޞ�\�[n����G�ɋ�mۻ�Ξ.���A7��`o�����
$8=E׸`���~��|b)�����iq���|<��L6],������yw6��O?�4@��w����W�2>9�f��s,"bby���������E��A4�0�C�����4��;����@`��	�
��s��������} ���;ktb��?�"h���Р.�"�Tljb�#��VK�F�s��н�#iw��BN&V��e؍��{J+�{��<X
p�z�5�'L~��mt�����_=7>�Ӷ��F<¢���[�	
C?����۷�Ѡc�NÿfǕ����Z-�Ev��J{{'��B?a e�ڢR2�A�T
����3�Y�D��-�A��z�_��K��Aώ���g��O��"i�칥�s-t4�^-c-�y����������m[.��@�l6�������~���d-l-�ֽ�٪�`�ԡ�vW %�OץA�����5��T:��ih�-����jc���)�utA��p���Zi6?u6��<W˅Z:��"��*���BG[Zolx��,�e��TK�n$�t�H)iP���J��?WK.ζ^k����֎Nُ-,����K�䩓'�V�ƨ3�l7��N6) �p�֌��N����;v�6_|�{v��6��щÿ�����O�6��/پm���TL�4
���&����w�|������O=���O��v��=�z��}���iTktX���0� ÑnԨ�t�Νt�Dn�ݶ��_�d�c;�D�������c����-b�&�8;2���"��3�<�?�쮻�X����_<�����{�W_�����o<��:���{�O�������vۧ���g�/c�[|�)����E<�_�֚�5jP]X����o~�7���uӚAHK��\�~}-?������JCcL����'�	t�5s����[�n��BA�e˩
�����yl��mBT+%�j<ciܕ�Wpc�Ʋ�$;P��`�O���r�L@��)�us[�����ta����@@���u��U&��։�?�E5K��`�,Ց��8q�f�)q0½���V ����W�ś6b]������Ǐ��-^�:K��ǌ�)]T��Rtx�JR����Ft?A�91|q���zp7��[�]�L�1�q��1,����v��JQ��zk��`���T��t.��)v���S]�'A�bm�J�tC��qx���zc`����9��U�L�c!<����+Ʀl(w�.�ںJ��;]I�3���+m�Ð������������~�|���� %���s�='���6��@�T�|~��k���tD:`��B~*��������l�����:2�C:���ZZst�E����	�F�����z�R,�-�`�������=����ַ��?���e���-�{ueE�T��
<�L�S�Jq���h�(�G����:��������ě�W^�ں���k۾�]�[�nM&�p�B�ׂ�Ka��� Ŀ���\wO�㦋�?p%!є�^}��`&p3�ͤ���B�{�[t�j���|���m-M�{Y�v�_�#j��4��[;:�N�nm��-:��c��>�л�C�J�j��L$�,	E*!���b�$	zP�h�b�Y`?��t��,+--���1���Ғ˶57V�\���[,"I%�IMuk��u{����YԨ�e�S�[��ή��0� K����Lgy��nQ!aLQ�0���y �;��+v��4i�Ƶ���⁳*]�EU5M���UO����E+W�mTKb�g3���A��3�s�`ي�c������%�#Ol�qvγOd=�R�X�h5ԜU3 ՎA9��וK�f�#pmv��\*ˉ���b^"h��{�k�1�p�2�^�C:�R�OY��f����ț	Iu$5)�r��,_܆���X\(��W_~�X�w��*"T?��ÿ���n��|��_z��ɬ�|�S�}�����,Z;� �-9���Ɛ�Tˤ��`����E7��MM��}Èa��&ɢe7�������a���{�b�_a3 �d�U{�ϡ'3�7���?��V�	"�q�f�����	P~��ß�ԧ����zy����VC��C�t�y��a�3]�,IP�۶m+��0!�|���8�*E���RI x��o�}��3��	TZ955ցvx���}V�4�~v��=����O�9��9��m��1��)<PY��@�Ȓ�}�j�"��s��$�kHP�AT���yk3]��ʶ�%U�2Î��>���O7� {OMMa9P���!�"I2G)PF܂�h���1f���L��050 �--t>#�l����ʕ+!��<����`.K7yF1�	5���6����X
�J�޽{��&�jA86�Ŝ���\��O	*���qNR�����S��k���מ�45��0)t��d��ԡ����u'��`&��c�e�dCCdSYv�6������+E@�T�:��_���1�Jk5�<�]��`v������!�婩D*�
��J�r�N�z�7�,���4���aM�F>;2�5S�M7���+נ�T���Zt��'��o~���. �x�߅��-��U.�*\��5�s�d(�ھW�V\�%n�DK�tr������H��a���K���tU�s�5QU'a�ә��S��]]�,�e�~��r~2�����8��o�p��m%ҩ ���T���R�������P���t��Sӡ���ޞ��@,X��(,�;A�YV\��~�de��#b�\�֮M�1y�=?
�5�$�S%z"���u>) ) lX��o�%Eq�x
�C��C}t���4�N��	I^w�;)Q;=��x�&ǵ���D�Ve�
X]U��M���~���˷����A��TD��B!�w�n
?X�{i3���С�J�����/�Ѓ������N �ӣ��1	^n���+���h^ͤ$!t�5�j����qC����g=��"�iN�������qʪs�n�T'	��;	�9_�+���4��W�е-��N&��Z��b6���c�܄�p����|���.(�6���� �0�g�KT���4�Zk:�jvɓl{��ȩW�d�K�dSo�21�4�.�y-��U%)FfKx-�BO��m1S�|!��͟�"I�B��C#����f`éCgkq���\tњeK��(9�Dx��������G��{c떷�.+��9v�������`3���W���~v������������@���mR,����
��:&�-��W�Б�*<`�`@���i�oq�$5�<�����*D���fp0�� F��x�:zF'6�U��"(<t�嗗���"��>���K/��p�́5�#O�N���{��>�ɛ�\,8::��OV�����7��"l�`Ж.Ǫ��P��X��T\�b��Ό�>�yt(q���c�͸�k���9$�!���J$��`ÄV≸�G�&�_�y|̓��� ������Nl-��Y�9s���7�*�6v��S�נ�l���>#IU�My��E?�Οu$D�Н.3y~�mx� C�[~B�k���E�)i��츰�񻫩�G��!��^����ր�f�9��1�Ə˄��ɜ9s�nl����X�	3Ϧ;�j�Ι/�c�\�"~ �#vR���[A�m�l��^��]J[ �1�����v�A���)����y�
V~f��-D�-����AV� 
�_�گu���iB?w�u��ŋ�Š�90�5#����@�ci"�5.V�I�J�����o-�6:�c��9C
�������3��:%� y��K�2�w 6���J��L�Ux�>��NMLfRtD�X.�s�|�XT%���d.�:<L\,���'YE����3�<ʏ���?Y��!��#vt%�9�j`���T �z���j'���Ѩ���r̪Z��K�`�`8�Ћ:6���i�S	�V)�9uzp)��
?vͪM��r��WvA�W�]��0
��>M�?��	!��L��*���z��.������fTt�1��c`��<�P�OgSZLv�Fg3%`Df�x�r�sLSsu��N���"!�|G�k5�g�Ux_�!yu8t5۱��Z�,`�L%c�C5 �*��	�"վ�خ�L�ѝ��v ��5�R��	S\|���IV���C~_�7bȁҦ��T�o����f���T���E�D"|d���'zu����wwv�0�u�Z�r�Z��9S+�^�kq�L�AWx��S�/�間����o�{�Ǌ����Jj-pN�R�%BDx���I��+��w��ִ$80��e(1�­��9Ӫ�q#�eԨ����?i�'֬Y�.�I��r�8Xr����CB�e4=S�_���Dl=�!���V-���\� �N�<(x���tA���	3�y��
�/P!E�d�� �|0?ZQ����F7*��~��cY�|ံ�j�:�|`Y���U��[�:�7؍�\Ĺ.J�W; ������G�d���[1)"$���$���1��0C136�^Д�K���bw��y���v�7Ys/�ӂ��ŏͳS������p-��p;�/ijj�t���U�� �������2a��ehF�s��L�"s���v���iR4��*�'�ܣ�\H>�s��P�}~������g�x����<����Ԧ���TU�E��Q<�!�| ;�����\�&���VH���w�0���-tww���rm��P�%e~K�"o:�۹�Fw`x}��8*nƸ��w ',?Y�CT�8!��n�Z*�G|��}�ʔ.,e�ѕsLG�T����)'�
S����^}���0M��N���qBjj,X���U����A:�/t��t����
8�:1��ǎ]v�e��l�z69p��ҥK�]c�O02�|�Bw���(����,�捫T��Gt�,�5�,ʊ{�+�N���	3n����JRjB���nIL�������:FR�dA1�9-6S��wu�/[��5J���>���f&����~�TNHL3��rͶ���sTx�--�dO���U��C-������g�kp)JS�1-����Ȯ׬w\�vA����o>��q�22~���E�sf2\(5�qv�b�>U�B�mG��+ϕ�9͎T�==}���֬Ϧs���N�X�����q@б��`�n�4Y�<f!?=Q+C�����)�����@u�̀��l���~Z���Pܖ)�
[H�{�:c.�u�
(��LUPΘ+����~x)��+"��ͶFc���/ϭ�Z���z�e+�jU���^��P��H��
CCC�\wG�r��D����RSb�
����<:G�u%Hc����D��4+���S=%�tE6T3O�S��bJ�hD
�nh���z��5�)-DRs��������i%T*>�W����زB���jI�<]r��r��48f��b��d*� ]��")�ƕb�a��}N�ȋ�h�)	a�h�|9e9h�HVA�Q�.�u�&�W�YdAS�������%]7-y��/b�]t��9��k���1��$5E�U�
Fp�đM�m��	����b�l�ֶ8%�wtSK�H��SW�)U,�1%۔a?$����w�M3ŏ}�����U�|�͙���lն�Uk��b(O�_(��91�[��94'���ɩ�'�V�j/\���?�y���/�߇�&�iS�~&�V�B����܎Ki�r��+�Y,�ĳt��eu�v�5)���d`��ǬZ)��7�H�@W�E ]p��@�ґ�jU�g��mͫW�����I7
�0�f���C�V!%���7n�͋��u��Λ�,r��O��� �����
i��w�p-�7��ѣGi�d��q��{�¬��Z�${��?S�&Gy�WUWuU�09HI����D����ɻ8�6^X68��^_�k�z�c��k�^��	�DFB	E�F����=���+��9g�{��Z=�U_}���=%�H�z���_�$�ꪫ�KS�R#��.W*+�K�#��
A���G`��hHz��t-�ҳ��2�2��-��6@W㻵:57�xƚ����~�z�H]��4�&� �_&�iZg���<�L�(�7P�a�U&�Q�\��u��*u���
N�`i#�|f�2��1���v$U+����.\X�l�N�����2(jٚOxg��������fE�BIx���%G�5�	˰7�C�>:YF�{뭷`Im��o��8�t��Y�ǆ{{{a%�v7|�W^y�СCk�t�Y�r��Ead)���OE���ÞM���;3�QH���)%��II#nu�5׀���.!pM��~۞=�<����;������3��'a��*�����Mu7�x�M�.�K�ղT�����.��^p����g����P��\�dJ��׿��n��;61F�C�\2ͱ`4���g����=��Vt��H�(.��ZGۜ'N]��V��ez�ZSS����13�;z��7�{+�>�h2���I�9���W�L��<�S��9�c�P}0�"�h_��g�~
�����zz{�������Lf�����\��Ԁ����4�J�ɩ�U�.���dy�'Qpk[s&;�OT��K�1Lq��r���'J�bks��&S��b9�}r�C���j%��l$e���?�ztll�e+�Lf�*��Q�e�Ю!�;e���4<ڔ&��j�2:4�tQ7^����h2.e�����=�zn*�G�&;	�c6a G���f�lj�@�L&����)\ķ`��������hڽ���~u�SUǮz45��c��?:>�b��s�/�^	��i��#~���3��������W��7�u߳�^�J���I�6��U7$�V	�Xle�z��R�z%#���QѠ66�Z^��x���㿹盔�D��o��&�}���=(����k��z��k׮}��/���/��?�6_�я�T7�`���ʹ�[n���a���XXS#��$�d������t�?��_����N.]ڝ�FU_�Us�߬˨J	�be�W��җ��]HEX�A�l�R�"7C}�`�M�_��C�x�{�9�fL�r4 �����+���Ts��ƛ��F��v�Õ�-����eȆY	�)�|��'_�X����F�J( X���)����C4!C�ϾO�~ɾ�d�&Dҟ3�~�
�k5HD<�U�&���G���w=yx��X����5�%�R|�g������S�y�c��
;�[ε��j%с�I|E:�i|���R���-�d�u.��?�tq,�q��@K�?��C��#P�����C�u��;#Y��T���$�[<v�(l���)�s�04!	iR�'��|x"ߟ���`5;��`��YX=�5;{���4��ܹs�Q���Γ�iii��v���$����Mb��R
�,��Q�m,��Z���<�Fғ
���>	Njg��8*ٷ����Ո@W,�䙞t<]p���#�} ����*T����+ǎ�.Y�����\�����_��Ȁ������>x����_��R"�*H���o}��K�)�r\�o�@�NNR�y��K��{�x���!O��#%�����@'�s�=-M��G�ߏ�_wݵ\�#m��o��f��%ج���P�r���fB�L�����R���v�|�'��ܷ����9Ϳ�ů_~a�׾��k���iMUJ�X�Rג��B�5%���`�qu�Z(㯟~�P�O��sN���o�p���q����O��X��A9������شiZ��\C"�f`�p���E��{>��������&)pi*��!mc�џ>}�-�J=_�%X�Νێ�����-��z�&�7(cdt�\���--@��
n��C���-oS��Lns���N�M5�m�::2~��	l{6���"�T�b��'����8�w�y�t]��(*�8CvAvblll�+ݰ{x�ys;'�G�N�����|T���1#��{w��s:�LO���,�X�b<+cv�(��h�PD���L��̙ɉ)�o�?	V/ˍ�M-��BQ7L�71<�s��5Q�
b4�N64��wσl���Bap��h�Dw��pC7�?��<"�τ����)�!!f�Zg�͊���-7������ M�#'��!��!�ܚ;^)���lQ�?}��P}Ƌ�n^{ٕ��qz�f�W�z�4Ba]�G@�$��وt��(��K�=��7��믿��];��P���C��_�r*�i��8r�4����w�(��٥��j1�B��/�Noߩ�\vŢ����Ç`��M���%XQ$DA42_��[o���'�2�z��\����P_���g?�����qˡၕ+W����rAFkl�`4��֭[�}�Y�j�_\{�J���C�x���� �>�6[�r�UxI��O�[H���޽x�
������o�P+��K��Ջ�;���(��XҙaP��.*�޷ou67`��;x��	���G?ʵ;�9s�����>}ZJL<͕�\����T���e��ch�!�/*j�j�� P8�	!���<[�.X�vh�s�l���T%v
y/1aB�G2E���}�Y��!�G�'�
���'��R,���4�/d�N�T�	�Tj�UT]�p1���N�(��z�6�V������ �HϊAlrqP���2}~xn����y�I>�!��f�u56RD]%XV+cO��ŷ�sj
�d�I��.�7[�2[&JINv� ���ݳӵ�`־)��h]tќ9�}/[����#5#�q�E)�3�1ʫ�>���#��߻����7\�kT(�3�w�� ��o������5>��7�x#j�����̓1�z�7��;��'7o���id�]���l�ʕ/�(S<��/Pƣ\1��ә���N�-[�P�߫��˖��mii�t`ρ���>2�+<��9T�~bH6�p�w�4��p��La�Tx��%���ckMԷ�Uȡ'������>�1H���;�钯Z�n!S�V�%�0�g��3�����5Q]i�e�OpE�BY�T����R�R�������cX�A��T���܉�S��G�&~V�(�R�Ec�&�����8�6h%c�t���r>;)�5խ;���4�R���!P
�yn"I?n͠���*����Nx�A�|(u/-�J,$%�|jA|��ʦ���:s#!B/�'�~;u�Z�DCA���z��/�x��H(4#Uc��иbϧyCR3W	��q|�T?��g �tṿ������@��S�sa,t��遐�z<�[�K.ܵ�h�!�f͚	����(;:�ҺU�z��P�C����t:�k����hz~Q�M�T�`8���u�:��ZE��l>���-,�lՀ����sfj�߱�XG�\����y�s/4�2��MdK���"zL�<~��[�})��A��{]B�����ּ���>�g:�΁g~�]wu͟_��
��Y��m��������n�j��kD����.^2��4R�R@�u˴İ-����K���)Ǝ�f�i%�G���kn�����/��N��#�e0�W�@	A�E���[�즜	��,�"Ex]J唆QQ�L9S���W����\�N�"�K8@��~��gcuŊR��=��3^��Y�x�
��l)O%�'N��>h�|65�$�"���8<�`����3�(	&Kl�Ƴ`�a�,B��A1qY�R��J�w"����bC�i�x����ɿR�{�H��:5[9�#$�
uv���R
��Dޤ�R��EVk�g�W8p
3[�OBĴ$��Ó��OSwgՋXhu%XJ=�>��X�� �����%Oم�I�{���O��7����}@1��l�Aa�x2�A]z&쐔���Ƒggh�Q����e*��UG�MB���@Μ' X��7�<ZLa���6�N5`%�=�nl�ڦx
9T����ok���-¹_z饥bt>��,"\f�F�2���z !Ѷ�аHIqz���$&2P�x�u�����D������.5�R��f�J�*���ئ={��ơHB�K^LAL�II8 ֮����]�j����*�o�1������=���-�s��
��*<Z��Z�I�C==�'ƨ�u۱]��M4v��njh��^�s��<+�"7������|"��غy�{���U+�UK�����GA��)O���4A�25������A�$��b�s��P�Ţ�Y&��YH�Z������s� �;���+F@�)P}SX���2B���R���C<�/���ʰF�)���ZV�k�"ov�p��ԭ4���zծsS?�l���q=�'�8ʰt��d�A�^�����/Mh@T*vͩI 	w�b�5Ŷ�!-�;Ye�:�Pkz2��N���J0��0WE���U�������'���#�{,�W,�a�`p��7u,[R5O<���c#���q�ƅ�W�Y�czI� /)���H �|�ʍ�X������ںـ� K�6|@�Ey4gP5JU�r�8�e������ ��F��H��u?3��]�J$���7$������+e>15�P8�|���o�}h���Tc�޽--M4�ϊ<��G��oӔ����::څ�px='O��b���V-�F�'���
���-_j	r$��11�%��"��<5����k?���2�vl�9���a�n޼Yb�l�:?<8�u� ��陚��;o��������|ʼ�s	�����'�?l"��.Z���"}�r�)�it,H~�PR�*�O7E����o=�|�#����6�OB�H��ϒi�<R�N��R��C�,�K-Q��,Q��?� �ѹ*�_����$�k4����
�0�����P�j�*�Ԁ��FHx����9�+�QI�7��[g3-:ښ�
d�uv�D�x��y�Y�p��N�;Gi糃�	�$�Yz�����Ii���2ГK�Xw�S���ș	mL��e[�M�-\��3%����ʤ����9�UX��!���S��x&�g_z�%��N�kE��L8���릹���r�*���ֈ������;��(#}��I���X &3�|�R���!6H�Q�NM�,=]_��[F�H�xѢ��N,��ēA�CCC~��\d4;��w�P�W�Y-EWn? �FcD�����v��1�������aÆy��Ȋ6�程��	���F�]s�L�.�<}�4np��^Xn�8C$��Q�	� ��B{z�C��	�DHߓ==��]�}��b)O�Hl�*v�B��v��J?���{�.�k4�:�JF��OTKŐR,Tt�iz�0dW'����>�_+>u���g&�둤Y���d�/[���il���T��-Ut?���`��Ij��&o���^�w�Z!?���ԫ�J=��\^��<t�I�)��D�m��+a	��R��H-aE6#-� 2����
�̠�b�b"z��U�x��Z9L�D��s/h"6�ʥ?T=J�)��z�]����V�
�AQ$T�s]�G�}l�)�?�C�T��h�j�8�V?
�m�&O,�jpώa�{5�e��,ؖ�����x&O�a2�aІ�w�������&�Vihi�����3�#c��|)��D�V�
M7wN�r۝�`U8�|���p�uqjh�ޑ܋!D#������5~����g�	+���t4W�㉸Ru*�&P�t@�֕���u|�P(���cP7,�#�F%����`͍1�����c�8�n��K�ݼ���ŋǆi�5׬�A��/^|��$(��}���}��>�s�0�'#��o~�켮{�G��`j�K�T��B��#+�-w�գ�&;"�\��pUq!���Iϯ1�?�ј���~Q��2�����ƑÍ.h�fKS+�BgG;OM:EVH�'g�Bq.V��X��Z�BH��dՅ3v<�������o��d�k`B�5$(K���\b���/���\��֩ZR)�SgF���u�]��_~�e,w���l��Bm�v�|���ښSb�A�y�xhb⋋%���?vp��]�;g����
C�Z��*�B�!��q��/g�{�Zf��IE8�M_��'An�b$?���X�Ak��;�P"���!aOi,��Lۮp�oP�i�:7�[l�Rړ�h��P\�[�ͮ
� �Sf�3<_f��JM
�$�G�8��}tFe�	���.{���7_�c]��B�Atxm<"*�B�8��iӦc�"�{e�0>�C���'>�`ԒjL�3�U�9��s�5��<g&7�t������S�8�N�8n��"Az��@��d_�:g�|���!�� s(�o�THa)I�����?���~���*h�����o_��װW\qEK[\zY��,���7�f�ѡa�}�PUh���ԤaX�p���������V*=��S`�P��+W��b�y�_���r���d�&�}��A��"	Z�d0;:�p�Z�r�7|��O.�w��ɷ�y��_���:��]%��r��f�g��&�Pnx$٘8��@~r��{n]��chr��ul3��Cw���e&��l��]�#C��]SK�,�V��RLH8���c�(�p5ujj�ن��?R2/Ε~v���98�Q�|�tpJ+39���x5Ű��(�\!VZ,[��9��K&�g�j���j9h��fSVT�� =<I�D�[}��^��2Y�s]�!ƤĴ$�å<w]��`����\�a:�%��$@��V꜂J�n�! "�Ʀ�)�.����.�j��㰏��iȌ]��ƭو�I�~����T���䦫����Tk�R�*9Z&G���ӓ�E�W,]�;�e˖T(�w��7v��>�׿�f�!3�Wsx��U�DX��[�w/ںo7�~��_�n]0�����eU�#1�D��C['<�b��niJWw���_��}q�՛�nz|d�ъ��}�}s�#.=#t}���~���W���_����C(�i�V������O~��<r�H{�e�6�gv��=�z>9����eQˤ�{3���Ӆ�kfsS��C͌L�<�W��Ca�V7<%�ük��x�����_7��L�"T�������1*Vq||˥���j�55�
 ��C�����\����N���{���S���w%�Q��ϋtN���c<j��k̟)2Y�y�w���;�c�?���2�yMS0�(�̸ђ�����\}S#p� �+uK�e?D���q�V���6�HE"�� ~���*�LR�v��AK��v˳_���F��x����#B+�*a�����$&	�&Ma�0���뜍�r��f���Ͳ�|�*-�R��\�kbn�6e
�xhx?_�1��"rG|i*�	Q&�㰆��Hj{Ƿ��ͮ�.r�c$ ��������w8� [��v��òpI�����
�n��Y�Z�Ap�@6���=x;(-���'sh?���D8p��֧?�i�=�/���8��'�,��V�i�x�	+���3Q��(���e2�D�U�o.��T�9�����O�[ߊYѻ��������ˎ�r��������ӟv�޽a�Ž'�{�_���5�"�[=��`j�<�o�>)$��V|]L8��*�hT��~�S<'(V��A&yp,fثS�u�blQeF67����ݟ��K.���t�y������4�[	�^cq�30J��'o[��#2JM���dc�Rt/>��Q�����]�~���o�Gu'��46����U��e�P�T��R�.;=�ڵx(M6��N(*�MՆ3�jT���l�*����g�l��G�v��Pі�x��i�z��fi�
��IgKE�_fc;I�[�J�G�L@գ�t�eE��8�C�ᠶ��X&q��Q��}9 ʋ�X͞��Qt�b�`""Ue��}#Ѵ����b9x��Upd`$Ю���,�~����h=��~���� �oѢ%�?���O@c@R���I�H�(��8-c�CЁZ��������|�37n,ש�����u�`(؟��RwC���L[3M�i�[��Sp�3��hC��jn)?�����voy��?ý���%���v~*㫚�:�R�HM��.g��T������o����3�
C�18�g���u���<��S�l�`]�X �T�����p�x���Dƛ��8>6�_�����084�޶�ÃC2J�1��LN}�S�z��/Z�+��LC��+�L&�����j(����=�L�g��fZ0P�e]|�?�~�C���7�Y�lх^����hr���P-8�f	$)�)�
Ǜ�Q`@��������p����u����r�-��]�O�!�^z��*ec����t͘E+�կ~EI��!ltr^7�;o��ꫯ��<��cS��!/��!����wh
Z�:�;H���M���!S �x�G[�y�U���M|�p8zο���o�M4h˕+��g"�2���FcR;*oJɈhfN��N���s��݋�j��r�M��PM���(DxC���le�xʯ`Dca~Q�ֱ���mx/�p�a��I�ָ~�G���=26�چ�p�x���Jy�'pAH���k_��T����y�رc�A�g5����d<�)�t��
^�ۿ�T�ŀ�	����n�_t�E���Y~t�q}N����g>���)�"t�(��(�����g�j�#	�
���\�`o���y7@�p�(t�vǚ[�k���6�龾�x��w�T˶�\�EH��a��پ���^|�����	z��/�sNg�m�s���J�3z����~�˟,]�t�����X��.�f]��WN�8��+����KQJ �P�uK3���z�q�d*�����}�.{8' &�o�:���V�qk�`�th%T�؆e�*�j��\e��t�
�����7�&����;��g��B5�(µ��tCs���U�x�����xK\��`��TlN�b9���%��s�r��ej|zrbzx����i������z^�áZ�ꪥ���I:J�q�b���ؤ4Ǧ��PbE�������r�L@ł]��UՈ%[��d�S�O�p��E�1��4��:h�H���Ni���JƦ�Uǋ'�٩:a3l�6b�NôcC�Ԫ�z&��Z��,4<88�/PO �}ꄒL�=e[�!$���}��zZј��թy���%X�lމ����B�ţ�P(��@B����J�6�kF�����e+���\~~���9*բ����[1=6U�-��4�^~����Q��istЍ�-�T�q��]O�5�1��-�	{O��j"ٌG910qb`k:A8H�� \���V�N|�=�^�-�W̴
,_}���:�kJ2�ȝ�dT�e��֦&ÝQ:vB@��h��U��b�"	��Sj!��#^(�Ö�z��(e!�Z����u����ݯ�@��
���0�B$�D.k�뙾��|��p����Ι�=66z�]wRV���2u���������=
��Mm�]��`�.�w���{����sϵ�^��<�|�X(��a)W���{�����Á�"n���r%�*��G�\
I��,�ʄSfS>5}�O$�!	��a��:KP�+��׿��x� �I����=l�z�Ė�R�%�CP�!H�'H{T��G���$A5��R̦(d��.�D���y����� X��|���u�g�zk���p�-+���7ކڿ���p�P!�֡CG >�>�i�u`ї_��r,��x��X��}4�J��9�&	Br����ϊe+�Tfy߉��W\N@�������4�P������
�����n2*,=h��k׍�ݻ����n��VX�8�B�@���t%��m�4�ť��/۸�y���Ǐ�d��w�ŗ\W!�sv ���`�Z�	��:L�8���аk��w�ۊ��b[�����-�|m��&� @0�'�W¼2�Y��@x1/L`3���MRj>Hq���1�����۷W+�7�|s|rF֓�{J*� j��1aZ��Ϝ��ܷ��v8dP��R��v��$��d(A�D0?�$p�[���s5Wg��JeDY�L4B�L�%W`������
k��g�}ɤ^D��yP�	�Z򐂧&�f����1�ܹ���`B�:4��g��W�¾�^�/@�
��$��Dgۋ�o��N��_	r q�Һ\"�KћJ��"X!
���{v�U���axB���k��|A���Rn� 
�]4�՜l~,�+F�{z)�$���r2�� =3�8�7�^XSꩀ���)_T�h�`a�Bv�♓�2Ù��%�RS�j�p�T߲�CQ�*��������v�m�d���IXM�������s���<���P�!k���������s���{bl���̼���+ �8K/I�Y�:��jP�������\�n1���(����3x�5��H��C��c�q#j�5L��Un_2V���!�t��閖ց��c�'��k�@����6mڼy3>���`����%X�fs{�j�n-���q�ݟ]s�J���s������9�+��<�)��@t&�U���]�1���r��eăv�������|��yE�&3�ذ{Ϯj������Bm��뮼<�3���ݒ�`agGG{n��x�\�$������ݠ(t@m��,GBd�����k��f|� ���"=Ԥ7�ZpǂJ�\�&�m�aՀU�����
��K��t͟O6?� z�\��˗�x��ߥ�,YƸ^1�/p��[�݋�f�?��koHwU*a��!7.4N�dÃ�4ToJN�R		F��RD�#o*H����\�#>��%�"ak�b�m|�.�R^��&���lK��P�2;�$*Ez ��^Z�dG	g%��P�|��e�����?���~
�j���N����se��KF������n�B��(��ئ���'�.Z	������/�����)jM��ol�/���^�ɉ̂���������w'<�T
�H��t����>�y\�)�7<� ����?������>�9�v�.[���Tώ;���E����1�&������"�����2E�u�)e�x�p΂��\��ٳ��O|���X�3Y��w܎+�o�`_A覲�X-������7Ş�\Z��|-@�P�d���M�]�����!j���0�&����y��{x���J�3�,Xq����}��᫮����^�;��.ƙgE!B��5(���݇g������L�\�}��w�فS��B��L��Q�@WW|�8�U�VP/�N@L'GH��({��gA	�%�9V��ʕ��pT�)v�_�@*�p/�yVҏ@�I����X��;�K�(�Yۓ*X]����ʮ?�N�P�V�33�\�H&�0�
���\vH&���0�W�C��y�O�\��Qp�e�М����Q�`�®	< ��*��|���.�,����G}�ϯ��/��?�ᦏ},�䠕��u���\�?Z��Ҧ��"�&<PXł���K�"�����3��"(��PK���941����̪U��|&&2o���#=pd��a����H�Vi+�ȩ���`�T�R2O��^���ɐz���6�tjϾ=`��EKeK�Wg��N��ά]s�d8�6���n�����֞���J~j*�l�y!+R)W�p�4��T2�!�L8`?�Ɗ����Jv��:�~0��`��ɨ�4}W��d�$M�h�=����V���y6�bzN���ݟnlnz��w�K�6\���+�l(�*c��AJ)MO�4�e�K�Hc�BQ=��=x��i���z�!�dX�H0���N��'�t��RBe�H@!�~p�pԈ����C�,������*Ԁ��/<����>[�^�x�� �?s����w�o�x[8���3��kz�O/�����}ϗ�%0獨Ej�(R㺍�i26\�X����@&��oB��湻M2b߁�ep:.O6��P�U��=����ɾ��n��@�:���>!Q/�*�rAnV#�ű{���DaJw�������R�*�%*z��% ��'6Vu��ko'���)�
x��+.��B�*�OƳ�t�M3۶mMo��*h!ݠ�����J엌%��mؔ^	H
��$��5���6qK;�������ι�3��aÆ��^5�=�G��XC�w�N�+��@��F��z ����N�I:�.�^j�K���n�����/S�a�d���"��f�j�,O���H�'�N����d��%�/2�W��ԝ�c_�D���xX����{�-��`0�ֽp)�B�����ll\{�Ň>8����'d��FF�(��(`���v�D��x =v������9 :>�s�@��I.l�&�G�E�K�����͍$��*��F�oU��;n]�z��%�P?��_�$|O`D�殮�]z��8�d��ԝ�e�5k�<�į�^_��!x�8�x��:Q�Ð:i����+�pM-(�Wj�d��ؔ�x��^�:(=�}�F�>�zwr�H�����XJ���2Gי��чS�8�I�o��#Q���0�G$N!�J�$#>g��s��!�j��Ć\(���
�֦VaW�c?$nד�t�B�kߩ<�H4�LE�yc���[��l�\�x�b�[������ۯ�|���}�Ը����nZ�C��tjѢnl��T��|b)?���d��0�3(�7��A
+W��f�j�~�e�(3UͰ���W�99Q��)���FD���Rx��e�U���H�=S��774RH?_�&P���-3���c�i���b����գ
o"����G����0��q�F0!�W�	D�S(@�� �q��t	�\�j�GLH�J�����B���������#3Pb|�s��jr�o�!*s}���n53A������j������IY�u/��hK����ѕ˗M�����r4N�I��Y.7��-���	�_7����Y4F�N�&�������k�F~���Ra&G3�R~�<�[����S���Q���%��9�s/�qϤʆ1�jAŭ��m�PWS`R[gGh�	Q#>��:\�@�����X�Aa6��D3�a�&��"z�]u��X��#������#?�J�tc(���j�,��LJ�ig_v�J"�[�^q�B0E��H��u��x�琪m���D"��:�y��@��� ���x<)U9WA�������%BV+��(�gy�z��|�ٯ�'&EX�ڵkS�4��O}w���of�����x+�_�ہ-��T������N66�۳���GB�Se �"��+����G^{�{?�) X�"~�8R�V���۱f8������+_��� �SZ�K|��d\� ���B!6D�����˯� �D2	�B��X�ě]���d���8\��jL�ڱc���$1�B�$T��:s�����Ƒ=Bĉ�ކ}3�$r$2��f����ረK� �|$`_���t�4��hd3b��[p)��'�jHP[��+4t�s�t���,�e�F�+U�����1�̒�B�@���)�"+���j��.46Y�������%� Я�-���_`�Tc�k�X�5i哩����}EJM���J=�p��X"ht"�i�j:m��m��&s��;�`AQ�&��x��1
�{a3��B1��u���T���}�!� �M�����E Y�qM���J��g?+�p<�{۶���������kZZ��G��T���/������LQ���"����i��f��T�����!nc5��x�>�AS������G�H������CM]p� ����[���CLLL�1ab14�,��i�ı�֖֮E����v8�/� �7.�:<ሔI8<pfP�)���qo��.]�,���������5�=�R�.l��0x����T#P�:��^��R��3Y��*���������B��Fܢ�c����%K]�f�����TҙN�9��[�f�#�1Y��5cgښ�O������T����R-�U��J\S�۔-f�t��P0l�akղI��~@�T�^�iZ�+���4n�/S�t��"����露*X��B�A#D]�PeoVJ��R*��Q��%��E8,�E~���Ȱ�w��|��L5��ɒ{���S��(�r۵S��Tzq�񊥊��s�C���
�F#q� �����%K�RǏ*���Ic�8e"O��L\�;Y��K �N-��'Ӎ��T�H� �	�
� >�gZ�m��`�n�)��,;�, (<f�_HZ$�:��$N�E2�p
a��q�፫ϰ�e,f+h���	~���?��?]x�J�,��{���O�3�i
���i>�8\�;߇�i����
��曗^z)��'7ڽ{4���?S��L�Ʀk.�����@�P;pV�9�g9q��֛�x�{si���7�]x~0 �L
���իW�\	U)U�̥�I���/;p�w�y���l�y ��iH|~�޽X�H���JB��3]��B|:�Hd�ҥ�3�>�"I��MT�����xG� ��\��~Q�H��d��T!0�XD<(�r3��þ*�D�o�\6�J�s�q`�W���˘ U�"�!t���k���#A9��!����ў+��1���x�k�y� E������%�ӱa�*�ܐ�I��c����X�"�o<o�$�'��@Z d�����%�B�'q_ɍ�0Cr��Y��㓠�P��|BA_�B-R�����X*JeAu~x���Ɂ�è 7ɑ�
�8�āj@�~�f6�b�d�c�`|<��2����,L��n��[o���H.�梵�POM��Ov�ݻ���V|�;߉+G�p�<6=��׃0"R���m�Z	!���6�2��2�& ���g��I�n�$�588��s��4�7���e$˼�N�]�,[^�|)�rj��h!&`�͝��o�`�|�%�0���L����`�\*��"�
�ʖN1\d��m���s��16454BS��Z��������'NصZ,� #B��gǚ�i
H����C�p�LX������������>|�EI_����!6�\S�k��b�H��1ͅ��% iP'�}��7u+����vO�ZѫW� � 43��G,s�YedB��ߩ/Ҡ�)��<|o6��
�r�.K�k��K!Ej��D��b�ʵrA��i�@������t���j�ftՅKN�=||ɒ�Q�T�[x~ϩߏ&N�A�=���F����I7�7,ڈ�D��A6���F�>.Oq0H�9Ĥt�b�H���wp ��]uU��,�OXsp4�P(�p�r�D��9��Skl$�i8�z>!�֔�ǧ�CӠ��Ѕݥ�����K�g;����눆��Mb<�%��F��p����c8'�)����_�;��я~$m4u��I"��}!����_A��z{��.��EȘ�4�	��4E{g[x4�9!q���Z�784�5HP$�#A`Q4j��֬Y�ZR��۪�t���9��YȤQp�
ںK�\(B<x��)%��M�I����#ř43I~R�������D��^�(�M��|�A�Ţ�~�9�Y������*�4BjH�)�]�"���ţ��ձ&*���4�HAF �(�e�Ylr��f�i���|#��b�Pu��oO&�+����~Su�C� *(JG�8��SI�69�*��L��!��d�n�a��0nj�,�8��!����BH��8V�੓�h>G<Q(eFr�P$��� ѰR�%Il�6���Ρ��%{.j_�e'��J��O��T~,bP�{͐~|�A����	���cs"^�Q-�#B�nie�B��2A��`?,�<Ћ1[	w��8;(�-���S���t�����hk��U��ٳ�p��:�r	Y�T*��-�����'�[�ۢ!��r������������أ@ݪZ�Z=%P��a��Rp�|I�9��l>'ы���-:�FV�5k\}�;��w��i�'p���J3��\�l1��?�K:�tӸt��!l���%F���>��Ҋ*s��e��ٮ�5��|�H<�����,����o�E�[ZZ���+��㉰P>���nI88iX�
Q>���hjT�j555��Q��Ǐ���As۷׸T>;3���R,�*6������J��D�]����r����S��#х]��q]�9ͦj1Xp�
��e#Ae��Tj.�E��� }���f���!V��\�q�M#`S�h���l���[�m�GU$�Պ�X���T���AU3�-���^]3�(Eʶǣ�)"%�Y�|�\/U_=r�;�}w`��9��b�)ݨM����O-�h���ޫ�n4�<�� �\�/7���h�J>u��Lb��手��;&��4�yr���☱]
�~�������m`�����T2�����$*��!&�ڶ4ȓ[�Ѐ/��.�����a�>)�A
��`{gǇ?���z^��#=0%�$œB���`��l�Z.GS����u�����(ή�?�������$���U/��:���z��Y�ʡT$�5@tA�w�s���V��ΖJ�B�}B�"=I�H{��ѧ�gĜ��~>�;yz� �=dz��2�W��M� �d�9<וW^)n � ����O}�S�A�ع�����uv���%Ӽ$_DSǹΐ��2�V#�Ӄǎ[�hv5�����˃��Ǐ�|�3���NOO�����:����(g�5S
g!��à�|{�e�A ���j|K�e<NCs������۷�>��]�W)\p�o��TSV��1���pM!���I)9�@A
ζ2r �?�4-�����ά|��B�9�#� �Vy)�0�B��]�tG�p��a8?v�|��u�P=gڈ����z�/���[v�̉^z�= �=��v�x�A8�bʉ�?��x�fF�0;��26:�z͚3���s���Q%�P�8;�_�j�Ny� ��;v���{{�������*Sa1����X����^s� ���m�����d�9u��>�����R�i�7�cH��]�3n���K����������������$��~f�T�TJ\[��8�hb��۷m�4^��*--�MsC�h,���L._��f���J�)�GA�ѹ�G"��Hl�Uz{{aoJ��:������ּ���Կ��`<�6��]�v]w���ց���x#b����L��*���7�	Ɔm�+��q���;8H�v�ԉ�K��{I��H(���g�X���D�Elo����7�<c���&l1c�BxP6���5�Ҁᩙݻw�.���΄)<:2䢨��>)�Ɯ����&@�A�cU�{�GF�lo���)��-���J��+;dJ�Z}K=�����Bִ-���.W~4 �,TK̄�]$9)� {�V�a�A��q|���OjN(bz�Ǧf��B�P*�~�R��
e����?4@�^�Y���E�b��!�MeřQ����{�����f*�@�R�S0a��n�ma����[J�YE���n���'��O�?�;?��SO=u`��d:����x��W��4����^�p�#�<!
�'�ɆޯV���9�s:n���_~�E�K��4�
�䩕a��O(Y�����?��OÝ��5�h��������/[K����h�S%��h,���~��V�#dE�,����?ݱc����T�ANH*�\\��*|	(^����$�[?�-���*)���y��5I���$� 
ƕŉ\P*��e�T�\�����)�^����52����'Àp�۶m�*�4pc1Wd�(rD��.Mi��@�34)�A��x|�b����_ܽ{�D���1�)�txܚ��:ؾ�:��Z[��;＃�b��Y�Vr����h���k�C�f �ʪ�+ث C��V��]l� �Ng[;�p��!�s�$�X'PIZ2���'�i���|E��@��֥l�c�������L(%V�:Ilq�t(Ȑs.Tr(��0���+�B�Y�㩳%�q�FV�~U
�����"Y�jL�gp�t�?�<�ӔVv�������)����'�`:h��ַ����r�-�ny�����^vrk)6�Y�M�6�t��k׮��n�*�J*N��T�v�ׂN~��'9(�����Tr��i���k�����_|��vu-�z�����n��'-�?=1��G��o��o>D�̌,]�d`h�f�#!��	�-��5�/۰������?<��������P�͜���M%5�_�u?kp|î�����#ƶs�H�V�dU���/��������[�a?}���>���)=T�lo&�P��;Z-ͭ��aO�±�T��c��d�z�$;��3���t2F��4SU�6h�H0Q-V�E&�FhR�o5� zICFM
4'�I�Ҕ UN�j�����a�����!Ai_ͩWaG9��
A^,p�C�+�P���	�J�ڛ����N��ի!͏��Jծz~��S-%`DB��$�����@�A=�-�8�d�������`5Ji�C)�U<I�7>ɍ���]vj���FxE�"��'s�r����5��Sc�0��T(��y�Zw�xm�����cajq����q�9G3t�V�;�#Շ�	Ԫ�T�UR
��4�x4Э��NEb�rɯQ
�u8�ѣQՆ��u��0�R�I��u�Tn��[�o�;ibv��x���xl\W�b�z�����i}\��Z���x:�-�Λ��*��]bW�Bi��o>��1���׾������ۛ��2&x�u�� ܷww�����>u�f�w��eW^���Q��zp�k~��;n�WO=����f5�+��k*a�1pXV�E]��s\�\2��̙�\f��ꫯ��ޱ�]�0�T�{t|Rlz
+�|�X���Źe ����@~�Yxa3҇)�VB�%v����R8_6�뮻�-[�n��={`2Awu�Ѭ<�i4
�CIm�����Q�j�F�rT��l&���;M��!�J�8�iK��U��S��I���)m��J��m �%�z.�F���P$����	Ռ�H��e�!��Sj�J��q�Ŝ�	����
+���+�?xA�I��SJtnx�������EO
.�Za�(�E�����h�\�V�s�yP��#��sY�[���@��	�H�x6��M!������	���U�%�B+�)H��"�S�2O��%�&#�i�H�����mY��$IFE�PtUE�P�S��~�X���3i2�P&IacA�۷��߸h^�F;���*LI@N��R�ԓN�S8`�?�Ǘ�ߵW�5�����o���?�1��ȑ#R�3��-�^�t���<�D6,J�@Zq�p�K�7".>y�7���{c��R�Fe��R�\d� ��r�Q:��hm��H$4-�Ϫ����@�z��x"\*�5���?v���F�n��C�����[oƽ9��=	}�/@�F�/�R�1�ܴ�;���]�3T�z�և���G���6�]��Ї/���Q��f�4#�rVQuӊԪu�%TA�%m�e���Jeo�'�$E�ε�yʨƣ4N�hzz&O�s����
��q���
��
��]���T�%b�C�(e&���Ve�)Ȁ `
v���ArJ�qI�^����J���'� �R;������5WL��e�+T�s��/��Y��{H7����C٫$($Y.�aO
S�r�e�p�B��.uHVŖ,�]#q4�6)��Bɣ�d=��I��ffJ���ⳉ���3��C�#��`@����J����A�fYTςd�ǊR�@�;��[�:��p�����5'��3���#��n�еw%�~�����HA�.����D[`���Y�LA
�uM�ڶm6����S�������}��}�;���?<�#e�I?X�����8��3gh~k(��舄^E�r�32\�c񚮘�ڗ_y���|��t(
q�KVD�� �'&"��珌KZ[[[�X ґ�V3��1�OJIw�!"��N������o�zg6���_�"T�=���7����|�'�QxÊ*��Q�ŒBg<ƢE�$��{�~͠��L��2�FM���T
Ez�� 5$�,�P��:�E1�蚈ҫ�hK*�7���wi�<W� ���|�RRW�?Ix�\�Г@?r��,�/�uW� Y�U��$~�G҅Ł�JE�K.N��$�$�V4���<�	�=����4�crM��]�L�⪉Q�Eq��W��z�As��hu9}i�p�I�y$�n��y�������p@x�R�}�w���~�c$fcU�*\w���(j!��B�RBŤ�Y0B�q�*RI���o�8l�rY���E��G`�-u�t'(�>� ��bE�M�[q���)���UZ=d�=W�Q"�p=�����~������֝PkC_��}����~n�v�����Ɖ�_���7���X��"�w��O����
w�ԗ/_��b	�P�ŭ{�Hxbl|NG�c��m�M�۷�x�U%�|��w�Zeͅ+3ى���T��j]��)�f1�$�'uF��w���{��~��߻��^�	�w�����찮�P6��u��B�2:6��lE�է�Ϗ�����o����涎O��ҹ"��X���@:��
�7�Ϲ>L&�Ǫ����G�p���X�
�	�-��rgf2�G�a�����p�i���
�T���$�%�zR��� �=�V���E�	�-�5��K6R�X�h�
�M�T�0K�ZVTp�eP8f�Q�^�+U���HA���b�����PY�g�q��$���cV�������(��Z�D����5Y�У����*��W�o��\��������_�D�Ɋ�"�:�Su�#�Z�?P5���2�\q=)抆In��Y8<1�	�.E��+Q;e$�ď����!ң�T���S��ԝ���͐?��J���x�dgU�Ě�BU+�i�U&�G)�j��	a�a���u����7�˫�8p �8|��K��{�Ƕl�K�O�sȅ|	��p�B��(��&�moi]�by"Q���H_����T�n�4�Jc2�H�i�n��㳳�@�u+V�~�͛7����r��ߩc5��^�:����@oH1G(L��P��U�dslm��mk%�y߾}_���O��v/^"Y���u��`3���<����E�rH8K�fݔ�[�a��M%%|���5\g:_#ͬ����-�"K��r�.(.�s�C�D���4v/W��UT�J<��K����5��,琍��0x��B���ϕ�H��~�ee'Д�m^[M��W"N�u�Q��8y�^�K�U)��X�(],�糵u��J9�(OQ�"\�r��_����T0ӑi�y`����A�FUaf/˖�^%!�гK���m�1⸎$��o/W�DSL�5��*���"T�ZxV�Q�U@s�|�X�$���0���J�#�M�����t��ڸqcGG�-B��Ԑ W D"��:�,����y��cǎ�v��59:��k�A<�\���;`,�ְ�������Q$-������=ݶ`���fJ�)\R�&�¹M�Ϊ��AJҲ�L�K�i"�]�FB�-[��2t�G��C-��	�;��9|�����Ujw2)@X:���>��ŗ���s�T���7m��b�s���������S��b�e嬱40pb����P��MF�N�>�������y�}��|f�|Ԫ�v/eZ!	�"�h"���^-G�m/�nn�)�����dL�~��8�8ٝ<u��ɓ�
���\\N��h��!U,T)rS���$� �Z|���*sj�� �!������
u�wK~vԙ�@aBs�a�V�,�1��+�{�c@;A�-�v
'De��ov��Pl�6,���L�$��.��϶�L}�'/����@)� �"f�BV}�2[pL�n77L�+ua��'%,T�����^R�9�J���U���PDi�"�V��YO�P��b[��zҧ�6���#�	l\ԥ�+��+Lf��|1��k�����cj�m��2<���"O5�11ׁ�	�͜�Q����63eϙ3����.�=�x����=z8kx��'�������� ��҅+W����3�YVr�p��a�6���������^`�\��.��f����`lc�26NB��-�
���ι�����S�p��#�Z���N~�{�G���GC�3��@��TO��;�'� ������f�����i�@�RK��a�O�Q�I��R~饗��ַ
����n��T����g	�i�
2�bO��e(J,Wk79v�[�26�h�ƍ�|zrj:�$ǭ�ފ/��|c�����Kp7:��ߚXL,Ɔ�^�x��:��"\�;��+v��53�*��k.>\N+9 y�f<��iP�Zi���lӦ��C�bqv�"�r�NP.юI��bxӳ3x޵����@O&�:�{���шȚ��Id(���Β6�V��1����
�s�lb�%L�-����@-��&UD9�d������j�b�$�[�6��Q �6Sx��PX�Tr�����$ �x�tq�U�� fP�p�#��T)R��m>-�F)ƃ(V��	zU�Ήp��r-R�s�G���}w�ȶ�2@ܟh$n��]�Ec4�o����D�PH����#G�`�3N�iq����p��B�i��E?����mE�[�������~���l���,��V�Z5=C�d�G��5�\�կ|����G���?n�ǮАXBh#�Ö��(�2�S��rm#��ʮ�}�O|�b������f�����.ʛ�Y��:'Z�4�f
'��R5��Rw\�Yo8�W���O��?F�s��Ï=q����<~��ߵ���K_�?����c���ЕX��V��M
����j9����=����?��"�~	��j(�R*��R+y��[���4���+���M�,�iTtT��8��be.�۾}{*LL>��.bM����h�J���8-�T�G��b����߰��Tw)������W�d���u�X-A�p�?�U�Z���t뉤	TZȚĞ�)r�ЈQ�|Nv��=�XXb28�\�|�}����L��M�7���gC�捦��:v9"3xJEP{\�X��/��K�,��<[vN�^���";[��R�d�pvZ��z������D`f���5ju	�="���q��z�Zmq*�Z�hU=�ɳ��8/��TT V�
BOr�k�D"�j���J53Ol�]c�z���^4<���7��4���e�gJ�tUW½ث*�	�Qثxp�'�#h�����Ʒ���޾���-7\���?�ѧ��3S33�0��v�$����~���5k�?222������K���]�7u��&��ۦ���{��Hlڸ���~B������E"����6��"��]�IUL�O�8qbrr���"J���E��p�;���w�m�q��{�R*,^�X�%P�$��g�tĞDyi��:<0|���ǦǊdT��]��6
1L.�����G3'*j�'&��4�yw��%K�g��ƓF��ށ�����rm��F�{��ԍ��]�l	nJ��-	��L�C1	�li�s���Z���dA�(I��͓��Uu�L�U�`#��K����ٜ�m��cq�q�ȿ�n�#Od@$�Ol48�ȅ�"D�wG�d[wH)	r֔Ύ�w�R�����:a�8�u&:iO���O���1	z�� @HcC�auJ�Bߢ�H��ZC�]���������B�V\o��`�&�NC53crmV�W�#�����O�-�������SF0�\��lcȂ0�E�ܽ�#�H,F�������~�ۇ[o�4��q���8�}���u�c�l��5��!�Q�!'��Y j�=p2֮]�np��55����������O���v�uÃ�� ����$ց�G^|�E��@�H��T��T��x�3��ps�<����}����]�ذ~�?�W�Ν۽{��N�W��x3_ ̗G��w�w���ի5��$�n���w��k_����=��H��
��s��X �c�ӧ'[�-���Ģ�x8�#̀uԃP��J���l؈G�)9Ͱm�VW������q���
1-�v�.��� �h����+6n�453E4J�+�I$�KN���/� !�;�� ���%ۅ�^�e�f�'��kp�����%IJҋ67'TTC˒߀�%!��P�s�R�\Ȗ4�������?[[�:R�U���B��8���qyކ��P�������q��1ړ�&sO�X('� +�����ȁd� ��Z��5[s3m.�R3�򘂡�?����R;_$�tNM�w*˧A��תN"�%�����[Ĺ�+�Ϭ��&�ߴ�Ԫ�7��MŲ�ժҹ�k���uO+W�����O��^d�_��W������ۺ�j�v�������j�:82��o�ʿ~�S����4`��qnە�i6�W㱮zs����?���9��B�jZ&s���	I0����S�^��w������7��ɋ%n��Wy䑓G��J��m�>V&�4��Y�q��ӧ��~�o�������5L���G�GG��o�R���8�O>����_��qE�3ǽ��0a�J�<vy��}�Y��(q�{����M�:�����6��ϛ�D
���{��OO]�~b"��8��D`�bŊ�+W���/�F�i 4E���	��Q}9M�˝�h�0N�&6G�D�CTQ�tE�t�7��)�I�'���dC��>�jg����ZK��j�x�H�%�R;w�HZ�l��;�����d�L� ��L��hi.8̥�HU�K�9N�$�+�4�U�
k5�V�"p��G:�~(!5g����~k��g<o��0��O�'�u�!���jO?�4=Z�9:����_z����H�����.3��
�C���#@`�(e8><9����K�͓��l��馛�ٱ#	��M*�b�vM�����,�5�&-ܡ�7�s�+�����:N-�F����q���lա���'"T칱�Ql�^x���D�y����f����\�|� ��&��ē��4W9�� �
��}������o~�ׯ]M� ~�����p���P	79���+291W,�+��n�b�".�fH*,SG��tj0M�I]y�S���V�ZJ4��\|�Z�Q55��'V�Z�H)����-��9x��O��ؐx8��Jy�zⰱ����)���L!�� 3Yᑱ{="��S"�i���L�,��h�+���Ǯ�%0+��^��%N��i��X�IR6�ՙ�����+r�Y�^��uXb��{�����i�Jn����9$p\�䭐i�T�X1D�n�r	�찫��Đ���<��B;��\0��9�,l��<�*@1�|[�
{�F�n�P� ��+	�U�R��Wf@07�I��n��T:7���HDˍ#FU�O�ʫ>���G~�-���a�Q�2�	��#�.
��F�<y��u�M7o-�
�/�f�+W�۽k��x�g>�_=�0!�b1	O�¥�c�؞;���k���2t|z�g������s��r=:��[Yp���f���G���o�e�|���fپ_������:U&�=�aJ���*b�"�?�:�i�I!;^U��Rm�f���:��R��ж����nlٲe{_~i�ƍ����"���l�~��Iiҡ��>m�8��͛��2��rL`+��ot����@��y��p��0��߿?�����~-��1�H`��X%�ʘ�q�AeL� o\�	�Ǆ� �x�t��6��Pk4���t��e�Ja�
W�ܭT�hk|0_Q����T,f"lR�XQ�2
�����G��p"z-�ۘ	'`22�֨J"G��	�͈V�%OA��0�����0	uJ,�
,�rD�o�,�n��A|i�gf	"�\�2^����,�,-��J���r���/��T�D��chS��hxȉdq�R�&�c|K�b���W�عs��O?62:����աv ��m�݆����"�a��Ku����'?��%�֒�U���������8s*E=���'�|��р���l�0/\�H��J�VãY?�F//`f����!���a���Y�g0��łvq2Y���M%��^j6����������q�"��X܇Ή���s�VJ!ޘ�)�x�ү~�k��N����+
�?��tW����̱�gn}ò��dva^W=��\>N�uv6�u�����I��<w��9p�!*� �Z��x�׭�>(-���k'���j��p��[c=�0����TY��#6��x��8�ڔ0�n?��L��Rgk�Xb�7���`� Е�U(���8uH2�SZ3���{� ��JH!��.ͩG�+�Y�x��	�R��d�)ٗd�=4ZM�pP���4�j�T��Me��m�w�ΙR3xF�`}�q�d4x�0����U�f�����IMx�ԍę�y(S�]`r:���t���Â�OU�D09�=>o��}��[n�%=y�^M�2�#��3'�8U�������O� \��=/0�Z$��J�G�BZ�,;(�d�~��q��Ɯ~���i��^$:O�����}�)j�Xmu���󶁭"��\�Q�[��
�uSLV�"���$��h�:g�d^�b\�RTi��Sӹ�,�����%FUh���ٶm[8N	�dW��{�c���Oo�!����BX*M���~;.K�j�#n6nO�<���TΜ9�1�Tөt ˊB���8f�������E���_�����W�-��I�%X�#���I)|�]��-�6��%��X�'�5n��&��f���i��I�L�f�Z+h�K���\� -���R)��J(���N�%u9r�Z�U�A(�$B(PL)�#�'2x��-3�k����ĸCzṷ��Z�q�2���|���ؓ�;d�uC�X'v�O�q�G0F�jg/L�D��Q�*�$��A0���}�#�6��v��ϟ�U�1�U*`�T�\�,�ENu\��2�N8�H5����&tT���H!�Gw�Z�*�Y��L^2�n[4�ϢA �&���4�r��9�ePsd��ґ����B,A�XRu�
�ί"D�2��Q����bn�~�6��syb.�WUj�y�Lm�d �RT��4���n�������qȨ,Y����?~���o�Ї>�.��5?k�{O�;w���~�SgvN�9�9uM�I!�����#`J��&/01����s�v�Yw�5q��ʕ"���p($���j==;o�0+W��}�*��T>9?�m_N�LN&�RU���r���.��i���+Q4�>��ٱl0����EF��Ǉ	R\����"	!w4�#��f��A�P�����V���(�U��Fg���
5�Ir��a��*:������=�q�m��('ah�qU�Dٕ�'9��F�!\��h܇\�@��'��Ԑ�()Uo2W4O�4��8�~+����\���@F�=B5�Z�^�[:�Kbk��Ҟj�aM1�F��1�h���ut�i��t���%��t�|a׌��r:�韝����ټ��e�ax��K�f��j�駟~���Ep���4�r�<�P/���+�Tͨr���Ѻ�i"h�b�(/iwV�� �?������R�����y|�O;HI���p�E�[i�k�CS�I�fl�8�:�}-�v�YG�vT${ͰM崞!�4�Jrd��M*"�� q�b��z�����I�fÆ�]v�⸅j�СC���wo�����f�C0<8^�����/��ۯ��k(0�a�>bC��ޤR5g�����'9�7���x������6A�^���0Y-6%��B�;�ta�L�Dwr�k�N�)\F������}f4�g���[���t��*7��<t�xj�Q�v��Q�]����,i�Ik��$�����B�*�DrH��R�$�8��
�Lk�$b���jIכiI+^	/��Aٚ-�A<4�O�+��m��]�n���BA�eb�/2�i�
٢:�#�\�TZV8j����?.�/	�:�k�%K�,߼��`�D�8�]��-+I��l���f��P�<�N��'��,
.��6H2�F� �~Q͖�$E�V����?/����$�9w<�\�2U9�(@�uG�� H'(�Sq�d���q~��G�%���dO6�����]����!�� ω�E �)S���j���U�T/R5vr��w��������[�4f{�����.�!��B�/5�=��O���ݣ ���Bgff�R}��M��~"7I�0�[�~.��E}��u�Nc��~q\�I�C���5*5�{�Q���Ȭ2�U>��ޑ�	��	8��:�H�t*
��	eh�)��%M��%G�F� J�;����;U�\!�_�/f{�$�v�:��\��R���´�/Z�-�EBp���4"�4l���0�v���aX4q�p0���D5%s�_Bl�%��E����w`�:������M4��SVd��Q�Q�p̨ԋV����eɛ����\��*xq5��h喭]<2�����L�N�K�0�����,a�$�C���@J�mJ�Y�P�����{��P=�*!�U>r]i�9s�F4�� �v�٧1a��/�g�A[ĐH�qt�pD ��p�PDS��� ;�cjce���띨7J���m�o�������
�Z��P�,�5��E[�Ǐ??1�dD���p/N2qa�Ϟ��eɈYIb�rL'!���9a�H���8�?Ecgw��
��Ħ@=�/^K~U�"ݼ��H:<�I��@�Pd˻���B��(����oiEs,Sl"��9�H�%X~K�@hŴ���9�j�ò��q�A�/��/)W��Y��wQޝ�Ǵv4���%���d�)r+�I��Q�6�FD�/Pl�x�"�"�8F��O�K�:me���E�UC�G>��$����JOT�
rm�n�9�aF�|� �O[�y�nV��I�Vu�:mll��.�a">�3E�ϣ���k׮ݿ�x�4-�~���Ymj�Xf��a8b�ĥ�O,���x����&ˋ�<������*D��!�d����`:���f�T�^�����S$��4����4l�����#��^�
����).�e�� P��P0^�\9����%1��s���|vf�8��z㍷*zN	��-�-{q.�������J��� th���j�\��%qA���7��1��;���� ]ިaAtC-W�cC�X��\��ϱ��i#$�C6X�ȟ�e9gæs�^�eV�5���UJ% í�����#`8a���xL`G�ѴD���IN���RԜ�:MB>�"N���fU��i��E,%�ؑ9��Az���	zF���<���JĈ�C@[�r�[l���=�����*2�����\��XW�K예"O55:lߚa�+�j'_��u�*Z�+;[�*�%QTPF�\�d__zͪ��C)�-�\���:��S���ԡ�+N}�kxfj���6����e���v5665&ާRP��G"!ס�,C�&�XG�ΗHL=@��pca3���z�ٰ�m�v�����P�4x4���L�$��L+ktq������59r��Db�´$¡ 	O�3�/,����U��;T�7���N�jJ4�,_���k�!��І���={ZǗ.]�iӦ+V@��Id�@�;�O&s�I{ٽr�t�K%�(�L���S�S(`q-�x5��Z���Ϡ��}�g�y_��tݽ)y��L��<lSB��]�#Ɩ�Er�\I��WNy�h���d���R]p>Y̬�gU��`Bjܢk��(�H:�-��� w����2w�rm��}8m�sIjܙ��\9?6I$��y�������Y��_��%���G��mY�'ԥD�l���cW��K0,������8z�(\�Բ�q�!k�+��H��.�4�9!@~Y�b���t�Nl��z�X��!������=݃�W\O:88�]�.�b8��t�������PBe�z��f���{-U+�s
5P�@@$�� 2��Tt��a��@��Jp#n������f���?��b�D���*�z�M����?nְ�J��푑���)#���޷n��'��b�)j��B�Z�D,��x�2��Tq8�}�`�RS��ny�B�V�{9����)�[�h��k �}ɱI[M>O���^��3v��	�熥4����i���d�i>��5�-^햄\��!�!�Ou�dU���Io�'a�+t=_U5��E6�M�L�)[��$�X�v���;��0I$�-�"X��5{���qy�(T'�Cm"	�y�=���Z��Or���	���2��?S��yp�g[#�^,F��Cv�iC��z�S�Tku)�r.��9A�`����Ҵ��!z
/%��Ö#���fs�fv�it�,�����L�����?ӵ�V���3sg'�ƾ���Q�a�Y���G}Wd�>�o�S�ȳ�
E�(�Dz�U�����q�����Da�(*1H}�47��t6���A��쨸%b
$_w��Rdߚ���&1h��K�)my�/�U�h�x�����+L�R-ep+b�W�3}�����ׄ�j'O�D�7:4
�z��Λ5�Hq���#G���f�/}���h0*�
N<N%<V��S�@�t���>�{zz���T:|2S��Q�B8�t�Ѝ �}-�,˔����1*�g8{a�|?��*׾Ĕ583I>��a6|0�"B%9	��6�Q�}��*OD��f�m�����������#�H��a H�
>�E���&b�V̑�V	�$�Q�Xbv��cC�³�`H�.�\���i�c{ˆ*�U�pH��I�B�0J�(Eӝv��j�!� iq=�)�N�Xy�VVU|
�S"I�V����;�4�]y����6����#���Z��z��߿�]�����=�lc]IY%�I�5FGG[�c_�x���*��@��L&�-��Hn���RY�MY.U3uB��84�q���7�|��j���$���~h���/����CՌ�~��m0@�l#X��Q��'NV�l��4u�H�]w�u�|��=��2)�kq�,��,��^{eϱP8����[�n�EZ˗.~��O<�a-P�9Uك��.�djzW�wpi�P"h�$�m��\�ΝS�E��l�7�����giڌ!����tWp�ـ3�.������.��2"ƛ�eA��r8���f���x���Z�h�ي2����n����S�F;],�U�.���mW��3��i��Lƣ\k��)�A�)LX��2|,��<�\|�f�!^��{��-P�'�KP��BM��@+���%6�p (��b��H�.�7�z:]&�_ɾȽ�+M������b�I�[v��xN�w���d���߈�%_Ćd�1�V����FKMm Q�����s�4�~pNݳ?3Л|GŲ���R�K�\����*2�4��o;u�u�l�[��Ɠ��=t��o{FSu8��|R�:z�P���A�qf�^��f�.R��0l���(��4X����4�4sa��D�'	
-��H�r=ŧ!�M�P4������;��9M��'f��J Kw�q����?�����C Aɡ)9���Q2O
�M�q�_��_�u�[q�	�!%fh�R8�kU�k����|���ϟ���+��5��()3G��� ��gF<�uQ
��C�u)�
İ���ƚV�
��ׯ������w�����ٜ���y���Ց� �֥�^zz��S�NU[5"	����mw�Sh����d������щ=l��S��N��r�GI.��n0>,(��f)��s�R�Y|Z��%��NR���o��CHh�WkL��o��(�Ԩ�J8�cno�?]�xZ����J4�ä���b
��>|\bW^��x���I:p�\GmJn���EzFQ�������J�N,���z��'&���ӓ��O���'�ܽ�xЇb֡C���i�kP�\�%vOO'���~����կ<r�v�Η_ݿo__� D�������w����-���ӓܷ��o{�>������,�F�n"L�<���p�^x��g�}V�gxR-J��7jx�k��L/�3�����?}��˖-{��}/������ir�1/�tS����;��/�"�P��@��(��a������m���~��������lۍ�_|���}�sمl}2���e��.<�pH%�I�4���k�⊹�8Gh��M����{����sKW������\v<��*�@�4�-8�#	Vå�.�b 5�s�γgOquJ*WTt[B'M4�xb&���[���l���R$�.�e.�S�.��O-���F�+I@s��x���%p������-! �ʜiur��!����à`��@�Ɯ\�T��I^G<7{inǟ�)���L�I:N���Q�3Νnl�E̚�CnZ�d�cq %�P��:�NQ$��u	eU���'�-֠F$Km�&5���}�Ő�������p�H�7�O���r��������"�^+:=w�_=��V!�=��ZZ�U��U>*���}��|�^���o���s/�������\�b���yж���r�/�瞿�����s�O?��cKW,�']i�ͫI��֬�dɒ�������p�̼[��˅�`_�V�N�"]����BTDd�l�B�5�oB��^�\��C9qͩy�
J��_���o|�@�p��C���/�%�)���@���M��@�5JK�4��:�V��Fh�����}�������'&pEF�p0x��������K��'D��tO�8�������=���>;K� �j�&�FW&Y8�رcX�h������U�VAѯY���0������^���zb�D�Q�7H	:W��]?(6P��F�Hi���Ō���֒�����7Qh�.�?*���,��CC�~���c,�g�XI�����Ir[v�x(R?��å���j��$	~+e	H5|���rWʘ"r1Y��i��'�#�B�嵺\�s������kyNF��J��x���0�{ j`JP1=d�|�՗.Y�$P�мM�ƫ��Np'P����u���tʋbe�]��Ȉ�iӦWw�ԧ>�ַݴ����^{�~��p(�b���Ϟx��������(�2x�[2w��=44��	�+����zw�k�ƍ�l�D�V���L6�?�U��TB��mܴ�[o� �e<��ŋ�]w����7ˍ�a��x�	l��d�Z-㥡,��5X+D�6��p�2�����k��v��!�RN��O$y���lC@��J��$��S���B�]#ɸ��Ϟ�h(s�����i>�`lfv�W/)\~�哓sj��G!�����k�JՀ-�iDց��Mgx���Z�n�������3' �F���2L�|z��5�;^�z9TF�V�#a�i����z����k.tVQ�7ʹk$x��K�a!G#6|�"�,����t��FQK�#n���7x;ƅɣ�\� �(d_h9�Y�����6(L�ڄ/䘶.�31��K�H�SbX��H4�t�F��&�?k�Ċ!�T���\�s���h�!�h�w'D>n#V=����=���]��&�\�Q�-|��I>c��|HɖJ4����m����R���N�r]��w�*g&g�׫F���E��ͨJ3w�'���I�c1�ի��﷾��Cȳn�%o�J�)�-ﳟ������l���Bnb�|��+����˃C���~</��|xx�ˮ%��z]ј62<������ו椩4#a�۴Q�U���+!�.NcO��=�$N���oU
�!mj�%�M$�c���s���/}��^�re_kࡇ~9;7�����_����2��l�4���+�B���J���_�pb��C��Ԧ��ޟ���wܱ��/�"@��`JV��r��["{]��Uh�bqK9;[��$�q�f����3#zڕ�b������3sP7C#���ƪ�"��iP���Ad�h7�l.�z7���=<��S*��/<��Kf���� ��Z��)U�����A�\��HD�_�>C�"�P"+� ���K���VA�I%�jSJK�(��&�P�嚟���.ߌd;%=&�W0.����o0�x�I��C���)x����b�MXΉ4ZC�5�a9�/���Rp��Yn���7�|݆�p�~�g؁���?���#����-��=|&)�����[o��z�5��T�7���}¿��W椺S8�����w��0Z�W���������~���3��$�4���l8Y8�� �X�������:,��]�LL^$��b9�>���[+�i�W>O6�*I{�Ax�aY/Y�������W�큔nؼ���^�|�|��_��?�=��3��Ξ??88h��>�к�%K��������	����%#�뮻����Xz��cbawXG �;�-�ҩ�S�x�e��_(��`���~��u��@��]=�$(�@�JU��dg�tE(��D3�L>'F�������R�Z����Z�J�������$*͖R�暰M-�
�Ei$�!���~��n�l��J���ag�m�Ht*@2GY���`�zS����Z%�0l�\�j-��C6�&6e'�/&��߳Ґ**���Xdm�CġC�m��b�&�Tx�	tlg��V��E�ZE�El$9,@|H�=�MȖ�ܩ'�m����.!�ܪ��R�*���tK��KeE�6�J=�{1��|f��'J��'�eVo۶�{�����km��A%�z����X,�ypM�97�n���|Ц�q������K.���#m�|���yF���4.�*�ӓL�#��<xp|bvÆM�#�4�<?���v���a1�B(�4e�uo8��⣏>Z���S�F�cz�ib��<��aE�~!3�O��я~�׶v�Zq��@��.\YB�n�����{����N��������M�å����5l��7�|�w>��%v�3$���p�J�QD��/qrb2��!��~;�ί�k��#˖e2^�.~��X�(��D.7JK ��0p�3�İ�C.dfp�Q��$yȍK��$M����(%Ήbf��'=�ֺ�^$q0�].nm5'�Tj厂���� �B�0/��5��z�÷��&��vߺ$�5U�t4nua~^�[9�E`%�n��S�HRr�xaIi]/�4ZMqV%Ym�=�0�vb��q��CB�J�d'����cy��q����b�D%�R�ْ�|�˃	�v{�4�w�L�
_4��'�8�,6o~㺫��� '�T,FۨJjC�E�2#�x��j��ҥKqB��o~�?����幹��W\����o���������'?	�a��𘤩���^�`_�8'�\<��^[M
�RN+���=��O�G�b�a��"�Q5/�U�+dҚۊG�V������U���#͒��ZQMF��q[�3�,�#�V��s�.��R��XW�ܹs�Ss>�����Z�n�⡡'�M,h�+�^YF4�T�|ڨU-(��XJ�|�������������l��?|�]7��b*�V5�,9�l�(d�X�h����l�
P֦��nl�m�R��2��g��уA;��֖
5%ǺL���=F�U�V%=��\/`qG$�OA�hU]�C&��:�⸽%�t�4��b�AQL=��)z��M�qO���j���c4��u��)D0�l�, b�+MGrӰ�)��+oenJ����q4���^+H��<�~\�A�?4��,�6��Q^��Sh,�R'\T$f"��C�N�J�D�.6W�T�ã��j9�f�}r���kB���vQu�ҋ���I#rH��TN��7��=6�7H�ߺ�#�&
c���!3�0lbZ(#%�����E���4���f�k�u%�#7��Sk�z��uɞ�څOШT-3��7Z��p]<ф+ՅT�őE����O���g3cc� B���:x�[�����;�;J�+�zZ�R���=���;��e�S{_y�F���bnt�/Q\�Q�3����u7�L�Ʊ�|D�a(���7� x��W���4jM��4�q.��@֗,Y�g��j��:�����<082H&�3T�23����	�㟓��)(�W_=I�RlĢ=8��/=�����"��u'�$q�%2�L�ഉ.E�c���[�m�J�vz.'���s\�C<�O���S:�7S�Z��!R7v�R�a2A�O	����ş����x��!����Ûk�IUH �¦ߔH�D���a��I�#&�.]'�SܹV�����RA�Ǌ8.�aA�֠%�����	��)|�T���+E ��b�	���E�=�e�&��N���,]E��<�O��|6r�$+c[��l�t*<))�[�j�����h�ZF3%��9sưm;�xCCC�	$ ���āԥ(Dp=f��|�7���л��nl������Ǐ�&�f�Z��������$u lW<)-8���+>v�Xxv
�<s�v�u�]y�:�e�,Jp�7����M�b�pZgO��Z�G�9;35>>
��
��(DΛ��_�q#܊..d�cc�3�bKA�/������R�4q����4c�=C�C�^z�%�;�I�\BI�����f�4jѱ�#�=��fg���Ջ/�]p֬�L�?���|�����ܺ�AI�ԒJS�tj��y����$�I�"�*)j�Q��Ƶ��u�f���j����ڹ3��[Q|�R��m1L�A���5XL�����LV��l��B��y&���d�
V�Q��?����D��7P.YMàu# ��WZ<��d0�0C�Pٝ��X9��L��$c�Z,R~Ҳ9�dR�.�+����ymn�N���nF���Ġ�٢<W�$�,I ���d�+��"�^�o��x%����>��	�������dx���t�ߋ�EU������b# ���U���=zu����}��khpz��C]-�T%�::�Jt�b����b�<:<zݵWc_|���|����s�n5��0:6&�,�t�'1??�O���Y��4���k������z�؉����J�:������:�ye��n�khR�
x����?�~�Mx�?��?߻w���'%	]h6�5ԥpg���@ϙQf���s��g>�b�p��a��_��_|��#Y��B��?�ѽ��+jR� ���XV#��͛���*�T`i�� �;w�\�h���2j��8s8O#R����.�S��P�;.�uf�V<K6�B��	ޜd���[h����^u�X�����zl?������Q�R��ł	:DN"�p�ݩ$�7����Iv�28��֦-��,9���c���$�8�8�����Wr?��܀X?�U�uR����Y���=wA�$�UK�A�t�Y�����6᷈� �b�(�'�$�w���d�bN-'i$J�Z����� �&z16�6�ӂ!Jq�P�Q�T��Ż�*v��=x19FS{m�v�ԅ7��n�n�}��W���O���H��?
�b0����"_�~}&��U=t�a�GG�'��2=z�(���-[��]|l���D\�{�'�|����L���V�V��8��}o�ʕk׮�)V�\N���
�L5��dx�;�����y�Qwh@.�7�?�яT����u�5[��5%ѕ������}�s���Z3�ـ#{�l��4�f�11~�Pnvpl�����/N�v���KW~��_֩���7����j�P,�ӝ"�]�a�/^p&���k�d_�Xl�x��N�˅���\����!B�ѩ��eoo�oi#ՈM�-I��D�B�S�Y�S�W�9WKS���1,
�EnhPJT�T�@(ac�s�E0(o���pר�T���Z�/'�Kƣ�=r������kSf1���rȭT5��>E���LeX�����?�jZf�n���q����$]��1wx��R����3oGR��G��3鍳�l��d2u�k4+�r�ɔ8��s�b1�(����,�B�A���!C�C�EƵ���c�Eq�-�V���	6Wk��VSW����ߺ�ȁ���Ӱ+�>DjN�/^�6��x�d��(�z�R��-��4�nv&�iӖÇ�����Φ�f6mڔ�gp�_��g���?�l�R,�袑�Ϟ�ݳ;>��O!����;��`?��z{�g��'��0��߫x�N�xw�����rj} w.�{m&�!<�׿��{�粫�Pe��������^z��ga���0~U����׮�����?nذ�7�ĭC�����}���!����"�� �xh�SG�}���?}vo���#���9h���X��,Z4��������^8x���/>��\�P$��M[�<)�L_�h!?#ښjY�ջ,�>#YY���$��Lp�	���U�a���BF,L�Y)��T���wK�2����%W��7h	�Ze��gH��x��=���%�g� )bݬ2�Y�	�mb+Q<� ���D���Wk�5v̑�m�2�;%���E���=!w�����^{.��Lu��m�܀*_q�=u�J���b��!�VrřżX,p|n�fwi�V'}�kW�ަ�D�xwx��[��;�G\{sxxWA���I^ٿ0==�dt�شU.�6{z��E8��up��D�?��R}^K��z{�4����� 3MJЁ}x�}��w���{�D�� 2��(���Q�E�Y�M�w/� &����7�Y��BwO?܊g�y�٪?q5���k���l�	B$v�ĉ�v<����e"z�vP�ٝMۚ������?���+�	N�>Mz�V_�|��_����^��?��O��{$��Vf=��x�����~���|��� ^F~���ɓ����#��W�"�KQ�x��Q#���ށ�d�;�l�X��Э��y�L'���(�m¼H8� �	�()e�սt�;�'�ٝ�A��!ك����dJ�:��,�+b�2�cJ�`ϳm`79�B�J���@(�w�Ar��č<B�cL��-�:0;�Z��(L9�Y5��t��Ĩ2ލ�#R����TG3�K_�y���Dc�	���j�c5��:��aCgӠ(�L��+"Ht�[��K���Z.��Pڄ��/	p{a_��d�\�*�䤎���Q<D�q�
�a}^���ߪU���xTT� >��p(V�C �ɱ���~�=q쬓�޸qc��?s�xoh=�VlQrb����\�Y�މGb4u[j+��u��1�U(���t3�O�O&d`����z�=�_�&w���K��Fu��[U�������ݻ���grv`ZR�=�"w��Wg"=j�ټe˱c��رctt���_8?	�:7u;�Va�@TH����i"R��n|880r�m7���Y�(aj(M�P�\r�%S�\&����|�&�W�h,�*dl˸�5�1'�Qg��O�I���`O��5�D\W".FO'r5-��i9�$�e��a��%e/~��ޟ��d�̎ږ.u�!��Lz��M{R�v����ŋ�~%��'����@<�8r��ǩU�0i�?E��� 1�4�k�u�=`�$={��#P��fº-�l���Z�H�+82��
�ҟ�n��zc�*a�H�,Z�Q��J3�bF>蹄�Re�~϶0�u
�%�$,�${��+妌��ӹ��2�c�p����[��S���)|v\Q��ݯ�

��[�uǩS�>�����^/3T(��#I�N�VB�x��d��c�M508̤[-}rrZ�:fs^�&^n*����������h�e"	�K	WqН<y�;y��W<���)1|�ΰ5٣L��=f��'&��1c��&am��=�!�	�aU1�؎���l�?�O�XR
��w���|bvǛo��>��o��~uppP�7
0�Q������'Y�r5��T;[�W?q�X����^@4����Ho�y�[�Z)�/6)��h��*Mxk�
#{�3e�"��B��%v �����NmC��j�r*�T_C%��J�BL ����B��l&M��A=hÞ�V�\���mRea��fpfO;Å����uvJ��*4t5_(	cR0Η��tlY����O�w��� �x�V�Gae���R��Kg��ߐ�8�qp�HXW�t=���pjq�=�(ת�8-r�\��DQ2�E�s�p��߸�D�Yx�w�kPU�L6RJQ۳���Q����"� j�H�e#�T2�*�Y`�X�1��*�?�v ���S�"!H�dD�M3*�l:������\�������u���/�әBE��Q�kl8E�u(�.3\{#�����<��Oɮ͛.�r�B�lzzѢQJ�|ČB��d��ASb�?���_}u/\�e˖Q��b�4�������]��^BFȡq�.ղ�����T��ҙ-*	n�[8�%������rA�3H.�%���a��Gm5ɳV4��5#t���'hvv�y钥��=����?�HE�7Σ��_��˾�W^����ccc��Gy���t�w����!�h5���%�[ş��8e3�Ň$���/1FNMM�ٔ>�r��O�Q�'у3�N�Blr��7I���l#ףɵ8��c(�[l6):�*P��P��M�F��b*���J���u��l�`ʄ)G�ѐ�T��pK�.������a�DwL��$4}�Ҋ0V��$���.qîl	�M*���O���tdRm[���ɲ
�EFi f$��:���a�`@1��H,�k��R�D�m�\.I�Q�����(R��G-4/k��7�	~YX�_e3H�>�c����}Y�(�aZq;��>�9O��%0��9�:X�s����d�!�صke�u�J4R��),_�<`�`�u��V8Q�W�eZ!(K@�Bojيnx.�SX�h�z%u�܌B�F���u�M���P4L��+LS4������ǻ-<�iȨqhm)�0=73�7\���,a���|�;1�j�_��Ggg_Ļ�/U���宙���H���Z�"��Πii����1��8�*"�X4��V�P�4�rV�Qo��S�a�|,���i�iWwO8/�KG5�q���X(P�7IU�����(^:�E�@u���J���&l]�n򐡘a�����硘V�^��w�5k��5������R�~�O�5�Ǳ�A�ù\oow(�89�m1���+Jx�DB�p��B��7���AS�!�q�`C��"<B>�`zJ���M&�K&��|	�:�
��E���xܯ߽%��{@i�����g�CG�h�!�z��O�B�!/hTl�����$W`�a4]	��4��R�z�7���LF@�LMO��^���I��"f�CX3+�������SG�둾��������¢x8ի���&"�S�^I�K�gnWw�U#�c ��Po�i��mҮ1��sM��CT�j�R�];�8?�`�R�l+�)�d/���UI��K.'��F�t���5�\�2v�	���8�N�Z��Ig$a�O\��0�G(P��i���v�|�U(��Jƕ�ٹ��>��{���L)���޿��/<��P����a۝={V&��M�tI�&�U$2�n1�׽nݺ��E�x�[�z��U[��/�L0:6��W��y!nضm����ʕ+��F����u�]c��<x���^�\�v-��e�^q��77xrF"A=���㩗/_��y��iX~I-^u�U6oiTk=����ۯ�f�+�y�ܹ��m�`<��_S����>��N�Ze=����/]������rV�;���x�6�ÿ~�߰\��v��c�ﰒؑ;w��u��s�+V�,���PϾo�>�~����������d�����g�y����KIu��.៘A�o��骔6���\6��c�M'%?�"9���4GM� On�Y�imvj��;�,'�}�*��Ti��
~]b
m�/����������O?}饗���5�\�s��4a7Y{�������e,�x(�u���4�ũ��w�8�b8L���ǈE��X1�Gy:_!;�٦3� ;�*IG�JH�ϋT��f�R}F���+i���QZ޵eG��H��M[W�g�2(��)����_�I�a{���m�LO�Ū9��l��1�H=��%ڀ-R���x_�3��Ą
�ŷl��Y�&���م\e.�˄"S3�o������ԺT�8�z�ݺg�ӕB1G�rfPХ�w�Z#ޕ���N�ЕW��pn�D,f�B�L�"��Db�d������4S!Ҫ�|2ٳj՚��E�gEB	���V,_���ۡ�T9����ٓ�Olذ��w��;q�$-�L
���a�ٛ<v��ǞشiӒ�+�=q��Yb���'��t�mX��_��ڵk�n�6�͏0qcoO<<�� ��`�-o��Zr{*5��a�f�9"|242�Z�l��]{`�V�Z�����;3~~tђn��j�XbѢE�'��U�!��+����=7;=��+t�ܝ��x3�du5��9m�mA�SD�C�۪�g���c����]"���@��RwaL���K;sҺU5�+�s��0~�%`�]-��vD	�bQ;b+�G��K�T��[rE�AR��։jl��ʊM�b&&���������a�%�5����Z���/�l{ټ�h��$�?L� |8�U����Zӳɭ����p?�Iɩ}��|LP��Y�w�警V�8��(�6�fC�Wŵ����02{���1C#E�f�P��� �V6'bE�5Aԡ�y�ۣ�d���=���J\#i_d�B�Ѫ�`��<5(��*�#N��ѣGc=h�U�Va������o���D(E��մ '��Qo�����;	c`L^x�7�i�����~�^��/���ϟ��~ a0ۄ�0����d`q�+��R`"���wS##�?�ĊV�-���+�>�,.:11	k�i��z�֭ǎCx�Q�p)q$l,'?��I�c����z���Pҳ�sx@�Y���m�Å�2�:t��~ M�������{�����>�����`����w�(Hoo���;~饗p����=����}�IDD�}�{��Da�ȃ�,r[�l�'�Uiޓ�/P$ɚ�[C'2f���B���*Ƿ����)��pu�?i�犋�+C����.�:�E�uC(�f�\��B���������A���&P�۶mWl���N8�+���&�RG�%;�k�^6D�D�%��x�R����RV�(�B��$���̀4�U�K~b�_P�X�$(������:n��49��٠)L�i�RKƘի�E�`>�!�)Z6�[7h�P�u����F��BEA���t�����2�����4�E��!�X��h�H;�bC�����~-��l'�r$��6j2���1�mt�^��Keh(��ӗRt�L��K��a�Km+���\z&�(��Zƺ�a�ۻw?D�\�T0L�={�R����u7'���ٞD��\*�t'b�0|�˖��Þf�~�7���3���򊫱	��9r��O|�^o�t�͹L��p �~�F K/��7  ��IDAT߸i3g����|wwO6K�2��a�N>�_�����m�$�4���`h�ϲ��F#�ߟ�,����k�V��ə��o۲�C��<���o~�3�BӁ��Zx��miw�y���8��K��Z�e����K�-����M.��j�%FV�٩
����3-�#�Q%WS�XF�*4�� �*Hm��mbW�5�'��C��\R�p���K`X�E�h&����������Z6_��߮���3�Ԑ�O��$����:Yb�]l�£���T�fB� �4�ӂ��ĪS�=]QiU��"v�H�(�=��lR�&�	�l��P"4F�X,\��cA�E�v�Lj.��7%�&:�JIL;�)2c�q�O�C��x��
���PK2ϖ�3HWִ��'���T�8����//�����gg�]ӒL��ڵk��5�~�{��l����+1�� K]Hq=aE�m޼�7I�Z�rB��I�nɧ	��H�Ȩ�A��NF�ז�dɒ7\{��O=������}p,�:�/�[�Ɩ�0X63�iǎ�N���F�m�F����
��{��Dq���o��޽{������/�H���e+W~���W�\!a�X-���+��� REt'� �[�/I[��]pN���oE#���i�ۭ���ۧ˨����Y��?�Mh-!�D5_T^��*U��)b&�Y�.EJ�iO��[�yvE�.$˦��,�A����Z)����y�]��V�VH�P�gA�߅l/N��okE�PF�������L,'�R5E����F���c	����r��r)��X��B|Qb+΍�b�
�%��P'3h3 ���g�Ƒ�[�e�۶gx�_S���T`b�p&�-�0_�}�" �U,�\�wm��N��F������n���fp@ ��
aD���������\K��k�:�dSuT�[.�w/	XAe~n�R��,Z��R��h,�Bjo"�>�p�Bl�D#���6�S�Vp
�b.Z6�����B��ӕjx�|%u�r�TP,�o���KO:7�S��-�=s�Q��F X�U���u��t��Q�.NL���|�w����7�9	W�+�$j�V:M��h2��/d����V(�zr�T�<�����+�O�~��?pv�����>�9�Ju_w��D2�h�_���S�T�����E˗\y�UpO�vb߾�W]q9��R*�%A����WJe,/�`n!Gm�v W��K�J��-ein3�Ii%z�ꭚ��/������֭^���v����n�i�ҥ;�|<7?���z�P.�-_Ȥ����k͔���� Wtx��'B�+��5
�=Ӆ�r,��0b�j43�r��':���.����Z�\Q[*y�&�ȵ�t�b�d�(DB4��Pi�jں�O�r.�ڪ랮h��鋰��٢��Z!B,̝�ļdSs��r%U�rh��7�5+������B+���T��[�7~�t��.�HӋ�S܍��7lL1��dI������͗��ې�Y��&!	�&!l!��4c��=.���"i��-��w��̗�<~������}O���i��<>��ԃ�)��q�<q�")���0�y|��X,L#�<U�a�@�T*�Q��t!�-��t{u7�v��i�6����P(�-��,+�7J��P�GU��Π]-O��J��T����z�F!�l>'5b�w:MuD�܅����z����b��բ�!�UgG������%��*d��O�X�Rz(�����?���u,+|B����C�C�㠬]�����`P/TʃS��{�Y*x��g5Ims}�4���?0&#l`�!T#��8��(X<���.���Ύ�_G<��z���w,��S!,����⊁��+����Ky��ɓ���֭�C�	��`�K_|�E<�M���wd�Ν0V�,� ~��7޸s�.�*BP\��;���2�/\OM�H�(J~�|R�۸q#����^��зVZR3DZ�*��B; >��,
��t��dͲ_���3Ss�A۵�ܴ�\�s�r�;%Ta(|Rj�t*����L�&a�BA����
p�\S����c����8�k^��+��@\����α���ؠt�\����io��j�(2���(�;�FH_��^ja� УV9éJ�����v:`����4¾ڔ,�lk�Jޏみ�������t�`�аu�(t�}^_�l֠8�ԣmفP�Y��+�0�x*�{lS D�4�mF�_!���̤�b�"DB�L��NG���U�)_��z=Tɉ�'�B���!"j0���NOF#�HW�YS��<�������=ՌA�cK4𥳐ooٛ��1Rf�j_�qk���0�>�����P��Bڮ�,�\>rb��}���w�^�h���˱�J�;3�^���[�喛�,��P}}=P��X�����KV�旿�?v��_�j">�撋#�u�<q��\���n�ʕ�r�C��RM��K�,���<~b�ҥ���#P/O9?86<2�����n}��K�[;�V����^��p���i���ǧ��������Y��X�񱑫�����611�u��뮹����#G���:���I��zzz�S),h ����\�yrj����'���V]x��w;~jB�U��J��LVO\�Ŋf����^�_e�9V��\L�+�Ӣ�<��0<�ȡ�+���Rl�mj��=j��@|<:Qj%��1��� 2%���2ͦ��"�]k�b�M�x���DU#���������%�����8o�N��ꋚ�VX���*&U��T�����W��(S�){vޛ�t�~0�;H��t��j���jghte��5v=�Nϴ6�am�e��e�0�U���Ux J�w:������޾�m۶uu�#McP����0b��{�C��˗
jA�$D��2��Ԛ*�����YD��Z��d� !�n�!n,� ���q.H��T;�۫�qݡ����8��a�H�G�@���6}�u��B:hT��	k�O'����B;.��¿��/����a�eКG�C$�g�8�9sj�ڵPQ�KXV,t�����[�����}� �}Ϟ=3I��9]4���W;v���	W�LN D△gϒ���"�ӜN6N<���߿꒵РG���h�5໨��!$;*�]hM,>�����I�9�w׮]������I~1"��<���S���/���o�ǡ�x@�O0�X�d2.���L�Pg�0�����A���h�!ä��pK��@,P�5K�/hLU�)Q��*��Vg�|琽LxC��"T���hjJ�lf+�𦒱jnl�I�5b�j�>~��i�����ra1}���� L��ܾ}{K5�X�2��t���R�J���dj�B�F���|���:!�uMM�JTp0�a�jH�g�O`�#�N|6���F�J�@�-���䧈7V�!���U؁��S/���o|���79M��*��Z[��{��?r�]w�h�&���	G ��rQ�� cѠ̺���6uA�+mD�e	I*��P �Ɏ�MLN���{����O�}7W⦞R�~�������%�J$r�"��.
FRp�u�Vw�Xʤ�x$�[������Ǐ�����&8Z�=���q���p� Մ�i�9zh��e��'r�̮�;��\���.r?l����}?��$ �2��Z��#By��7%�������p���@ȋ@���~1���������7�G���:�G���I���Ή'���I���|�wަ\b�r��~<��cGZZ[��ߋ/��O�8�{���[���z�wu�=}�ȡP����s�����ԀgL&�S3	�h<E�����3Je��lj湧��"�z��ċ/<��5��4��\(և#��r���bS�&��jN|i�b�%��5���m�d�|�ɓ����+³h\n��E�l��zJ���0��jb�ũ�ub�BYT�� �e��'�E*�9Ye��җ��e�z�l�Y4�]��c建B�����]����S%��8��;�Ⱦ��ϛ����V^�80x�Rm�ΤR��pCMKihj��"h����ǦϾ���{���vs�4L��?��wo���p=��@�v��MMN�:�uX�b��W^=��긭m1�u��^}�嗏ݝK��:;x$�Q�574:�S��
�PV6��������L&�y睑�C��t�����w��,�+���ƙ����ԴpT���������W���o���v��U�H���!��>���>��]�탒FJ��QF�5b!.�?3C��	��7,¹	(��O�+R�i˱z�j)%�<^�����yJ��4M�b��Lͻ�$2�)��5�%S-;�PNU�hl������,PC�=�+uj˰,a�)�`�g
�q�Flm�y������z�w��X��&��0x�,� b1�ӕL�~8��|�а҂�]��𼂓�3
4VEF)˓R�H����Ә2��J�	o+��!$�-ƍZ�"�\��H��a��$�*����*�vV��f� A�Hg��dU& ��ީZ�ڰ�R�Ps����G��G���B�OLB%R��"1��7����+�Dl����[,�_�z�:0�����8�8A�6¸á�����2�z����!��Uǚ5k~���[��VM8�}��~ �R���׾v�G>H�b��Vc���#�h��[o���������~�3�yR΢��)&��L��Kgr����/�ᡤa�pt$�z?rx�}�6]��ݽ�=r(����mX�L:e����w^`Oxbt�_y�����?����~K*��2��W�v�G>J��R�ه�ȳ%��b:-�	�!JOO�OF����NI�*��7���O�����L qx!~0�NU�MxO�J��3w�V�&(��x}��a�.'ϑ'@OLY�2����b>�LZ����a��B1�P71:ƽE��o���
Tu��4��� �T!���*X�l��ȩ
"l��pO��ؠb���b�M�4��<A�R"%�i�l�V���^���C��K�����4U�J�$�z[�P-r�.B{���P�;�1"?��4aD�X�M�Ag�7,��Md N��$MH�4�ǀ!��̠0�4�ψ���b�z����ĸc<J����kA��E9gE�k��0gi�m��Y �x����Jd2#�E��t͗�6��
J�?��=�~����O�Br�,�D#�Y�1��U�>w~:�q�<4�����)a74��̵
c -��3���o���߾馛o�v�?��Ž��>x=�����'AO����3%B�}����_�����ڦ�i�Jcs�(#��y��8o?y������jC���K�[�ܮ�$*(�P���;�Dp��q�yՊap��@v�����ttrɒ%8�XDl�|8��*�%Ü�H���<�<�:�����BU��.�@z�U���`:�RI�
���M����Vq��,잏o�җ���ۿ��������7�<zqΌ��RQf'��CpRT��|һ()S6��o�Z�iF0R�"�� �D���0J�Ɔ�id��i��2|�Q�ǣ^��޿9N��Tp�T(�|W�����:'w�2&�JeI!���9|��C�����H6V�r�d�v���.kB�X�d$�&��Ie<	�#P��J���:�o�FKz�8�!P��R8\y������
䲪�#�) �)ۙ�f�n%3��n\t���z��h2+�*P���)L��u�ޞ^���\�j�e�]�9iLX�u����Z=��(�X₹"�J��Y��F������{��^xj��yI�<�̳w�}�L��Z���B�ǆ�9R���x�ɉ��<�e�1C<��@+/Z�y����P�DI����*��y�_u��]{�ǏÊ�X�b�+��-͍�m�0�B��pc���:�G�ԼA.���=���.���O}���ֶ|�s��"T���������:�ϝ�M�����.|�F�m����F
�ݾ��ݻM�H��`��;�?�Ń��*q���%��>Ty$�M����FmT*�袄�$�x��d��K�\�
'�]4����R�}^q�**%�5"1Q\\˩2���%p�$]��	P>�ȶ�ǳ%�T.���g���j�W�P��w`���R�ޑ�2ے+� ��cʳoݳMCf�(�!��ϴ��LH�^���1���/>9>�-�!n�"Xp�T�v&��d��W�[�II:��T�G�ŤA0�N�t�U�o����qm�+��Q�ฎs��Xe\wkBWIF��)<:)�r��M-�{�@�р�R~��L��,��
٠!���Ln���JS]xAr2[�����|g���lO�/�~/�8^>�5�2VC|"ZJ��Sa`�G$ n'\6K���UM5ޢD0�[bj�8a���<��L>|��0�ǎ���:�s���6]�WUU"��LW<._br*��t��=��K/�;��d�~��ʬgM
��3�	� ����-��˥K��c�!����!�{���<��_��'?��}߹����� g��g��C����å�>�P�!-��?��kn����a^ʦ�����__u����߰i����6��A�<4L�_Uf���RhR��ѥ�If�Py�O}��J�����&���T�r{(�1��^9]v�Z���nMf0PP�
�q�\����\S���%����l�Q�Cb��YaI6R�5�Gm�	�a�u֖͚Qn�,���e��r0��S�;"�"#)�g(��Pi��/e��m���R�ĿC�0�\2��G��A�UU��&�2��T��0����m�Q�Rd#f1ʄ�Й?�-�2��*�^��Ρ8�@Q�Ql��d>�8P�/F�?�A&X�*m�Q+��F~���-��h�&���އ½��ĶCn������ӱ�X!_���~�y��K.����V�^�����Xq�EX�Tj��[nA��3��p��P!n�^�ڀ�.^�������_�~�GFFF ��������\n����tģQ����nll­/\�_O&[�ژ�*�[���N�<�Ȃ%�?��Of3�7�؁���=��{�7�/�3��9	e
q�]	���'~xh��9l�3Y���;}��.ްw��_?x`Aߝo,���(,f౤���)��bɠ1o�Y(��ǥ���i��t>���8�) �ς��rd��s�8)��κ�8\5�	*kW��̋��.��U�0�L���.��3D��wR�'�Z�d�<�M�%����(��U������C�J���<�BWT��Z1k���KٝdۥJ[�Z]���q����Li�)Ec�%� 54�D�CC�y@K�m��~��QU򅒋`R�!
1�HS�"����:�dr���΅R�Tq8��Np0G�x0 �KC3t����"B���Cq�F���n:���4Wy�X���,�'3��fX#�@���y5g4�51�}����Vy�����5��bX�+W]�x��jޣm%f`�>��쫲q��������s����~�����_������ڵk�x≭[�?zg�z�e~�jSC�i�
b�iM�����̂N?� �\1K�;�\��'�9{��
�<<|\2�ا�f�4�_���O�G�
�{|�l�<00�JN�R���u�mEm�u��կ>���ؿ��a����?�ч���,o�`�\"������f��+�`�i��i�l|�;�<5s���˯!AC�*�?��0����Zԡ�HA�UA
Y����M���!!+<vȡզU�;ʄ�bd�<�"'��V�`q%���.gCU#e!��RIt��6IV�Qdr'�'����β3�uH�Y��mb��$
��1˙-�̵;���E_M���d�K� U�|rr\J|���N&��8ߤ)��M#�����B---xVcR�.wV�_$.�t��H���8�B5�j�t�l76�I�Ǳ������/_���E)��`��h�f���^E���L�t9wI��I@�aQ|�ɓ'�B3[U�A��ֈê"�44
p<ϧ�{�[���u���zw��?�����o��?��K.׀݊dwww�F��BR������Ŋ�2##�mmM�mђ�sL����B�!n�U�����6�d3��t.[��СC=�PsS|���18r�H��6py�VU����XU;�.�u��~�c���n�g_|�Y�s"A��˗S�j!_�r�'-�0�J��������H##)������l>��˙�����c/?5�[��_��o�7�)W:A)}j� )�ԹD�e�.	Y���X�n�����K�f1,�ܔ�u��ݤz�SQ�E18� �u�U;_,�YGx�B0\��[A!n�2�(q���"9 ,�Ba31��V�kߤL�6�Lh�HV)��	���LGr��p��C���5 �%2�W����P;!������/����Յ�rppP36�t�

1�D�J���Q��H^���T�����u��{`M��Ӕ�2l�agG+�Z���4�v�|��2>Ls���%T���6��p?�'|U�O���Ԍ��q$�B����.e	��M?�Y��Q�A��u�	v2�Z��
�������W��z=������)�_U�D��r����u�-A�9� 0���eˈ�}o6K����s2��Y�d�������w��W/_�D|uxK�B.�J�@�.�P��������SG�^P��خ������H8JN�U&�I~'�J�c�d�2�.O&��'hC��s�>/�G2�����R�K�l�����ġH�H��k��f��o|�_�������̓���W�ր?L�����W�7o�����D�
����˸+�Ooo/>��[o�X|��G�1839:>q�`%(ѠZ�X�!",��޲yW�f���u������+�q���b̹�2�5���$��Bs$�E�u�
��b��K�B�`b�ɳr����8�W��Uй2}�s����Sҝ�)PW�o�Ó"�e袷qɴjW$�JмB��i8E�K/���ku���K/]w���c[� ��BEcup|��K'�>+v�W^�Ih�5\z饽�|�@j2����P��-[� �����'����۽y�f�D�җ^|z�����;���̣���p��|��>�52�E��O� �{}�u��%(��?>��6E�Z�(ע_ҕ��!5٤Si��C�Tƛ�X`	�� ���R`����X;i4���"��S�
�*Ư������֊U��������1����W����G��^I
�q�8@4��$��(�j<�?x��[���9vu��vqm�#@9 �A��0������|s��K���}�Fx��͍�|�������҄T��/�$�#�GU��f���c����yw������w~d�s�=��~WD�Ef�TI�W �>U>��N�I�T��3�{�cc=}�+W�l�_�0F�o�j	v����E�Ȥa�Z�$m٬V���`Z���g�,M����br5*��U!��}�
�#��٤Gsh�.C�`mpm�J/��w<s��q�D%X����ҿ�$lN!�R��ő%L���&�T�zR�$��c��6V#�Τ��P$Il(<a�"+Y��2RZ�Z,P�����`���q�LB�2v-���*��ca��J5[(⹓�T�������p��H~_ 86Fj7V3���𸱒TLV�GNa$(���+Vtvv=z�<����By]��7m|����p��ڣ������G�H$�Fơp���%V��|r�)}�*�WLNcP�'���<�u�4���T-�ӛ�EJ��T2W���x�\2���܉�y�{(y�Ӕ��������C�?s�g�Ϸ�7|%�r�m�ｻ��o^�l�e��ܴL���ؿ�m��[�l����DK���M�[����J^QTM���.JL*Z��4�;8'��?��k֯��@�Ij�ң�>
y����t�"�g�ރ�Op����I��3�Q0��画�n���>�{��?��/��rĐp¨���N�u�i���'>9S�Z�d����v�_�뮻���Lg)��Ƴ5J�`P�	�h��Oy8�+�3JB��b0�����z��(S�%l���L%�S�ԛ�?B>�piB�-��򹍀B�@ (0&w�r�S����K]*5�$i_$Oԡ��sB��d��l9����<�%5NӋ�-3���K�o㻥J`c=u{TL*fHJS�+b��8��;Y7A��0���e� 681�����=x��E 	�+�������e���A�o�8�wӎ�`$5�M�걘Ę�������t�������b/ur��A�T���oj�s_�3��"Ԭ�7�<IF�h�.G_�U4Ԅ9;�R�ZBWQ��,n�.\��o~3�x�>���-[6oټ������_��Hd�._(�g�y^dwOO2I�I�ԩ�8�Ј��Z�����e�yn`` ��Ą������%����8�����;�h�������^��|%L���nY������V������Q���P��$�#���y�m������}&XW�)�����~������E�]Z1+���Of�話��>z#FE��
9����r����޽���P.~"�u���	���i�5��hS[o����~q��|��J64z.�uE`�Y�l��% ||^�^<N���I�E����d
_����]��u�.!�)�%?�J���q?�Y�R�G('�Cy<�'W��A%aÅjգ<ڥ�*V@�i�dg+�T��v9=�<'%].�X�`5ݥU���21�Yf���j�*|�,��R�ɀU�;ۆ�����a`s����&M��r������A�!����&���az�:C<� ��|.�Gwh�M��̩��bQJ��:/��ʫ>�ߘ+L�TC���L�������4u���d�u�R����V��^��L�p�uk7^���a%��#�Ə|�6a��KV&�-d�M�w�v���8z�s����ʦ�:se� ���U%4��Zݺ���L��n4�6�^��b~�﷞|�_S�Aw̪U8W0C���փ�rUq�v�TʦZ,C�}����ϼ|�M7��W������|2�����p3���^��_�`����������G?�=��#��{��s��>��A�o������1�;��H�Pc���U�U��1��	���
���o�2�E��[$Q��F�K��|�M8��-���9ů�B�����������!B]BP�q*?��ô�� \#('�҈�`ww7^G(�@y^�vP�>\�����/}�K��{n>z�h}}�iyhq��ao(��É���cF*�xlMe_�1��غ(`A��N��[�J^���p��QX/�R��9��a��X�l���C �#�塺H���\��t��R^�I�o��U�K�tB[���UԢIĄ��-�)Y{A��&H1����)Sx�ߪ�.Q�r�8I�F�bL�>,l=��QDxa��� aU-�~�5k.߰aC<A���bJ��)v	���`�/�)B����C�N�tm�r뭷�
g���s�ܙ��]�J?V_/�꧟~��_������>�:~��,?���Ĝ�ʕ.�WR�"�!�6
��L�<�'Vpp05��7����9�c{�L��������ݻwW:T����2���:Jf^*�e{�1˿~�[��,�(H.�D��ϱzR���4=0�}���b�pzzM�Q���E�'q����_~q��}�֭��-��p����{��y�/��:���kl��i��C'��\&������O"�������r�������b�5�>v�(6x�]C��X�����N��<��?�.�G��R�e�Rd��ܟ:��1r�x<~�N���@63���}A8���A�q��Lz4W(�G(ÑM���6TQ5m1e��fTjn�TqZ�Q��GN���c�*��DD�zg�LR~���'��:4:�e���V	��V�i�b�d�0C:�2,��
���|<�����u�U���C��I��g�O�`h:�n--���ɼ�lL�\*+�z��`�ς�<����p�f�dN#l1���&��p ���u�@sQ�!�3Fp�,S��FEQ��M�3I:Eo��%Y����G��N%g�)â�U��I$'&�b�0�e��L5�l����.aE<�x��@�744�鄹�'��8��;e����s�*�#=��͖�@����W��_;��t{{{ߖ���ү�Νi����r��r[���RIb^e����wcA֬Y��7�8?~����trυEزey�������կ}۶m���D#S�<J��x4��8z��g�}���N���F�[�l�Rh�a3dƅ���򗿼��Km�� xł����� z����H\
4]�K/��ҳ/�n(���Tqi�7�$̠�IP�h}3��H�'$��j%�8��bxٹʛ(������5��49�Rax����`7���@��ܭ�M��ƳYL�hPPl��LB�W�I�2+�B-�Ҋ!�A��G��բ�����H��(I�q��Fg�<oP6�LB����$<�-�V_��%�IV�D�R	ةX6~k�2��RpeM������Z�Y+u�J.Wp��e�3Wut�(2RR��4>����*��3'���~pYAl����ǩ&�-�p�I�t���Уq����NN�tL!��in똏�6G��Х#��/Yf}fRIIJ�X��ӟ���84uX��~JˈT�4��eC�_y@YX3p#�cU���{]��wl8q�����Ou]i�RF=n Ȯ�/� ^g�A�t�׾��5+V]s�5{�9�k׮��~ٲe�md�q�_ ;X���#p���׭�t�ƍ����[2J���������;�����u	j��hN]C kW-��v��L�y���
�u_!��jG(d�uw��tܶ+G����"��R�F�BOO����7��5M�ix�]�)]�%F��LF��dL��	�TȗΟ�\���y7�:��"+g�n5W9��"�j>?���t=<>1�t��F!���fS8u�H6�q�G��Gf������쐏"+��t�â���5]ĉ$4zN�ǆ�f����%�%�������P8�a�U��%�!��f���kK�a؟�8T&�k$Q"x@5��1,�J%�0����n��J����<��%���?h�,��%Y9��aR�fE5lCp3OZ�)N��_�d��ŋ���ut�G�Ν;���8�8.U�,y"9�ĩ5�J���%�{��H0��9x�ܹ�W��h�Jn�"��֩���;^z����U�.�����MOM���B莦�8op��uR)B��ݳ�|��Q�\�\w��S�3Wb%�%�k:Ķ1�YL��?< 4�NM���
*�b�����=��)BU��ˣy$ʐČ�u,x���G���>�VZ!�u��*�mŒh1
d,�����,�����o���/@����j#:��AD��D��I�=����X21��6kR	�I! #�d��7'qB����3�HT:�<c`��M|k< ��( F��@%�d���p�����u�a��g�?n�
�XŕO�ɇ�"EA��Co��e���/���WC�>���?��n)��#e��<�@�e�R�9K��2t!'I�Ed�J�ij�Y��ikie�-���H�.�V�~��h��ڸAN����ò�Ȫ����/U�,����҂W��	|/�"����%0���jL�D�̣Q
�ݬB����x��˴b�����������Ƅ
Z�󸃡 @j�չ��!A. ���.X{�R��L�����S����ڢ���:X6���;9s���G�47,ϴ",~٠�O�<iVif�����J�.30�~�j8��@2�ԙ�x7�-��ŋ�h�I(S�"U�ǍSs0FJs�-
�ʠ�[���\��83 �Y,�l��|�\��K���@���鰕K�Ip(��O
�$���!�*l8�$����'�&�{���=�f��̼Eg#�Qg��y
t��s(9ꬷ-f W�g���ƨ�V	8�+�
���g�Cηa��|D E�7���,����m,�0�jծ�F����>� u�C]��MC ��#"M��ޠ�yhF�й�w����.��.B�����_޻��BQ]�����7T�<=��$���O;�{�b��+�pSѥj�
��L:��c��;�3r~ ��CM�-"�����s�	m�e�뛎'.�tݹ�!9-�ccc���b09qO�<�O�k��N��5g�m?\O�|)�/�E}a4������+�8�+/Xq����!
���D28:�hN>���4v�3��I�u���ZcM ~�RZ�HMn��(��B � �[��$"uq�&.�U�ӵ.��҅z�x���>6ì��d
*��s^ 萂��T&7��]4���R� ЉH7�/D���P�,Q]vu�\���XC";v���T[�ġL�gA���.H@[��t/����}�� �d���BK^��@�;Wԑ�Y����{�a�M�ٵĹqkW�a�`h+����a���)��rO�Lr���`�&�dW,����&[���3y*#yU�q�u��t�J��*>���L�	?Tv*���iښS�+UG���EÈ�wI[C����ӫ2E�x���%��S<��4$t�1 
7�q)�ഄ�u��VJ�2�i��Pz��?D�t>4�a�>�e؂T��'>q��͊��s�)9��{�������W�����O3��
t�s�YjgUnL�;D�ThX��~���BN&�p�(M�?��S�8޳��{��v���\#E��Gn�㣏��k��w�w�~&_*B���-�������<�����o��g� ����M�6�
������M7����?��ꫯ^���'�����c\y����Ss��)�lժU����Q�E¿x�bH~GG'dOȹe��;�I,>+k(���5&�ܐ��j��ʓ<$z�袋pZf��*�gT��#A�9������y���w�}W����R��̟?�֭�H=���O�6e&������~���+�wpA,VxϞ�0&���Z?bX�=���۰���a2Ξ=��?>�����tI�v���˸��,g�Vc=͋U�^`���,g=��S�LA�����{���%�Tu8j�F��"i8���fg�,�^=��^ۋ��m�������zj�Ũ�\J̥P%_2�1���� ��d�����`��i&����+QUb�������
�\;x�0:�J���LO@�V�O<�����+/g>��;֯���]n��%����EFI�O��l��<u���{>q/���oO��+[[ꗔ͗+J�X$o��+���:��P�~o��P��:�"сs���O��������GihD���z�5[�#��=��_�b������^��~wSS�֭�nܸ	¶c�[8m��qg*?r�t��[?`���f8�����D<'
�+���������S����䂾E_��ױJ������Up��Ϝz/DGG��gR�����2Ed�:q��%����.�
����:�Q�������6���|�J!�^4J�\�If�;#�N�	�'�,����!b��A ���H�R����B�e���N���O��A��r<�4��S2.V�2�l��0mt>�� A)۬Ӕ�D������y��G~�w��p�S��������=P'����b��U��CM�'�ߺ(f�H�J�|61d�&=��@�R=?95<���0n������7(+�3�7?	�M��$��
�K�ؒ�KSSX�s�R�y�⢝���ӛ�`�H�R5d8�FӿU�6=5�E���-�Z)U�~��R-�W��&YI(=�GM�kTc�+���(�Vq0�Ce�a
g�i��5+�νL� ?pN��3�{�s�\Us'��;%}'�F�T*��R-nomXN'��nl���w���)v>S`
���*�J�  A��qt^z��_�l)���}���ᘞ�{��e3'��믿��m۶����n1�~����objR����'p
�'D)x'�F�d���cǎ�"�*¢	c;�PA����uo���8��_"�ܤ<��C�E�w��B�v(x\7�c�{������Qڿ�X*�!�l�$i�ܩ U�ow�L�P�J,X��/��X�
x�P�b}$ܢA�#�^Ƞo�*ކ�L7_G1���S���3M A��$u_Ln�P��|jt�6:�I?Ciꀧ�P�	k��+$�2@�r������;wn��;���n��R�!��^�bH߬R�L�H�WFK���|�����G�����Mj���b� ���B��5�/9��.}�s��5�8
N�E�4��ӵ�YAM�:�W��M!�5�����Za"]���w#LML"�A�u"��7LG�6n2�N;4��X&���T�ȴs��ū�Rmš�SS8^�V��sg�''.����+.W��g�t��R�\U��Bip�ESA�m�=n�϶>E`��E�v�`#�w�\�| �i�ő�������l)m866�e�殞��'O������E��ãX��O���S!�*j���������OM�o���'�������F���w�y�-W�5ݱc;Dh��k~�a��W�8ߋ�.�=�'NЉ�zΝ��38?��1*%�cǎ�k�\�jաC�dvt�Òb���#����3�	q�p;��;��TOQCE5ʖ��0�j:2 OdddHXE��f��%�<6>�z��d:KE�l&
�?pݍ��e�_����	�����Q2Jm틱��5��XK���o��i>�.x��t6���U�}���D6��R���G4*^h�fofif%Uu��0�c���@���46B}$�E�#�k�\�:b������r� ��ֵG�)��pOy!��Q�"�g���F|�>rؤ���$��$��rɔz�E�"=�5���Fc��*Zg�F����v+�b�F���\&i�Qm.��̎zBn�*6cY��u�4b���}q2;A�W���<	�����jr���F)UM�ޤ��#ҍ'�B����41f�QV�����$��@L� F��V�$��n�lظ|`` �z����<r��=ƎJY/��3 !��#���O��B���u�Y���Y�
��$i�C:?p}�I7�p�(��_��_ʭ�����>�)�'��?�a(�7�|���3TՄ{��P���fX�&Y��	���/B&aۡ�qoB�!�;>�P
w++o٦��w	�tw@v
������!�'N�z"�����:�"2/ٙ�_~9��wJU)�_�����p�UB(������+8aXl^��Y���հ�;w���O�bMx^"כ�Y�ӭ��^�k_�$x��ǜ���OɰR2���4�V�Z.@dF�S�7�A�e�C��6�S�.>�:�11�L5��,GE�J��$���O'V��ef�H��
�r5���]KDC$?���,�;�E��a�Ee0D�o]N�S�vk:і)��C'��$L1�u�rE8E
Y?D�F� �����SuX�磛.�H[� _"D�z��,L1>N���H��Kp�Lc�*ٚR5JP�tqN���t(9?q��.(�m[��np��횮Z�����шm��-�e��{�0��B�*[�,�~�ݝ��|i���s��݅�].󺺝��P2�.=���u������?_�p1By��;2<���MR�s���` %-�w\�l��R�P��T�����7�>���|��%�Ǐ�DP����������p�y��\�l�:�z�?��+.���d���}���?�鲫 �D�T�>L�!	JJ�GH�itς�P8�����Ӊa%F�^��K1��=�ĵ��nio��h�?},���C-ݡln2�8{~���ЭD�C�>9,l&MlX�����8��?� �����xܪ���i���>F�̵!I��IC�pjav��\��#�l��eZ�$<h�Y�y���g�%D�6�7��8��'�@#���Xcsf�mE]��+p�T�!c��\.U���~U)� 2B�ʔ*W�56M��2#[	}�ۛ���R��	M��4�x*�%��t�T�%Ө�GCY�\,Q��r @��"�;��E ��	�YK�"8C�N��T�Ʒ�_�7�r��9�XC�DSl!=�R��-T	ył���t&+U2q�$3&�8�u��x��w�w.Y��
	��}�v�V������^0��$5I;���Ԕ�e*��K��8{��?���������xR�o�>��櫶,_q���#�1e�N����U��pD��xv|>.n>���+�@\q��.X� _==5��Z �>�bŊp]tpp���1���?�/��/��pdw�`]~��@2J�e[�r��F%�0|ݩ3gcm�#������04T�T�pC���	��ȃY�%��h���aU�p�. ^����;�rxF,ֿ��+�(��/Lĉ;ϥy�x��g��f*6��qH�r?v�i��W�\�H$����%xZ*��C��X1�P�X4ܿ���b5�Wnimĺ��I[�=ȳ�`6p�_�#��\ �y�IN��͗��}��U�l)�|�%���U��r�_��f�9�E*��.h�W(��)\8����o0X��~	]� Z��h#���3x�?�R��<*�O�W��>�$g�&���иM-d%1|��J�
�SÉ�ڕ�a��ʪ����F�zV�l:-Y���0~�E�s�ң�Ȧҥi[)����������C�W�fN�3SSu�mɑ�Yu����._�TZ���Ě�\�FI|�������ݻw|tԫ�'''�x�o�Ƿ�~��=�Μ:'j||ҡP)\b}8���6�2�̟?��Ͼ����~¶o߁�W]������BN�ԩLj��u���"�c��d>�߸a��g�zN,~�h�R�=��?{�̦-[�����خ�%�MM�&8q��A��a��&'��gϞ��f�P&���m�ڵ؅����EqI�*,U�u�o���ʎX�m�$W*<�cͥ����=y�x)���MMC�I۔��ۓ�e'��g�-^����U��Tp�2������o~��>1�D<�(4)(�&�0YXh��A%���vl"mI��S�ݽ�/�g��	��w8,(��^߁��W�Yfn�[�����2�D��?x,���������-������>s��o��:-��p�h�$��f@%	���)	�,Q��a�˭!�c�S�SԼ�xVh B���25<�O�����%v�f��	��i��G5��J�A �ɎJ<J��ʍ7�x�W6E$�u|o��������͛7�P�F�<���N�uKX-(�
� �Ș<��{����uMs���Fq:4bu�d}^B�H����{��Q\�x�k/������/��NB�vt� ��xUB����UVu08mp�pd���.�U�a9M�����a�h?EG� �46G8
�҃��Y���D�!Fz���K.��_���ç����;�q��K.�_�����>��>{�4�:�� 5��������[�!�n �)�:�/i;w�����̙7�J�i��t�	NH��d5�� �7*Hڝ���qx�$�U�	�Uĭ$��J�#py��0A�=����9m��O�Lx���q4�4�OR�x�믿�O��F8a�6T�#�<B�'M}Ă"��XH(����G��xC;;�qA�f2�)�]�yeժ"v[(�*ܺ���rږ���ڵ�s.��G�$�E�ĉ�6h�s�w�f�aU$X��)>Ֆ�S�9毧�|:-�"n�	�����Q璪��K���M��>}����0�T�$:*�r]����p�M�"�P��tO�g
V����-7݌�����}���u��۰aCsc˾���y����{�3���ǣ#�?�я:[�F�gsi��w~,��:��O~����$��*ݗv�N��n�4WK3�����	�)ei;��V�"�yS�s�@������ug�ld���MO���u"�IL�Y��ԑ#�U����ޫhzb*��o�3��	K���S�S	X�l}����[݊�t3q�Ӥ�bt�k��g?].��Hikk:xp��Ço����W-��[ ���������i�e���y
fΡ+E�:���׮[��O�R3���dxp����8�۶m[�����5����Rl����Ϩ��Ke�I:�U"�t��t��8�J�f����n�|3��]����r���+U�]Q�K�:s3���\�R&W�Ϥ�Ã-��rQ�$���g�N�'W-�Z�pd�9	n���>��,���	z"!D�Q۴:����}�X��q�nO&����3�b������ĳNg��j�2jN̄Cz*SX�jQ{W�ׯ�
�"��\>ĉ���ʖ\��eh~o��K�r¼��ºr�S��`Hq�<J�q�� ������[+d�az�ԣo�\�r����R��;�z��KX�Ww�4��%+�C|��%�<�cӷa�F��r����QjD�����KI}���>�۾��/��)U�Z�Ѧ����6���i��K�e��d#���A$f�g�����oH/T+VY+���Ky }�)�3uv�	�~��Ǎ����Dq�=v�kǎ#C�x'�:E�4k�lȐ�믿��w�t%���'�o-\��ߥ6�_��#\=�4���4��.���H���';gXSSS���G!�+:k��-A�мy|�I1��p��p���Q��E5Y��T��\�?�x.M]����E��3����\*�������9r�Hj&+�q�t�H=pK��&&�Xz*As[a��~�iӢ` �9n���� x��C��@�a����K��3�<C�hT2i���`E~�a��	T�pQ�! xw,��(=����+�k����>�����@f�(i�Z���ڐ	^1&t F�d}clӦMۻe�ÓO>�+cm-fd����A���4{�Gv���u/b��n�����{���m�ܺu�ukG�·�~�%Fzb���C.�9�����C2��t��#0�\�ǽ����gq��܈U�
�C�W<��ljҥ^��z��Wt�r�շ�nx�Œ	�UU��a�$m唊�gFQE3���Ą�.!�K�#�n��(N7D}��M8��C#6�8�R(?�U}/��b��w��(v5�ԓ�p��7/ZҀM��Ǟ���Z�291p�G���8�pA��ޯ|6ׯ+�mJM��innn�s�f|b�g�m�%ܭ���'O��)���~����~g˦�_��℄�屗p;�V�7�§ �a"e���bz=~쫇��+�7�Y���4��x�(��m�}�R������t�[&�"���ɧ9'�iin����4.Ϻڑ�G!�Dd�����9W*��0�cȉ4��Eh>��cH��2�$90~�ո����'S)�+j.�.�i���P�����f��2UL`�
�B��0�y����h,��Z����H��'|���1qS1)���P��i �� �(��V���A�7�MW,���9�u��ӡ��˖ (=��6_�y��bQ�044H�n��Z[Z[����%�C�z�{_v��X�����bj{���3�Q,���  *����8E�O��,���}N
�	z�0iA�H���?`4��0U����R�r-�B@�px(�P��'4�2�Tgg�3��P��"�#o����ᇧE3	���D
*?�7m���6��i���$N�7TU5<:u,�L<n�k�ٲe��8#�#/��|"Q��.�^�U���.��Ώ̛���
��gs#�٫I
[Rdm���}�ݢ��W�\yᲥ���g�]b�������UW]����g�Ln��88>VUh�իW߰m۳}��%Ĕ���+(��M	���b�&(�
JF�b��4�;��qz�6Ep�5k�������=<jǼ��?�T�i�P��j|�!�5P��z�[�2�H�;|t�B��2Y(=��A1w]����_�O�|�N���� �o���������ӸL�-뎏C%��b)#5R"2e��-�L�ӹ�����F�3�
�����ʪ��X���0����"G�XD	�(������z�R�����6����i*WlBfy��1�~y�[����Po,NU�4p��u8.� Ős����+�ǩ��qs�� b�e��&NR�`�Y��O0�|&�o�A"�I�W�)8�-�J��pOR��d��F^�M�rU!t��?��������B�0�4>�'[�w�y��eˊ��x���>8&��K�Xi���W3��C�И�Pi���=���uzЏm����N8�m�%���;�h�ja�^9�~"��S��������KwN����omo���(�b�I�=��]�ea�C���0�U �	ДX�֖f�/D������W��C�K��,��{���w�����+�O�v;S���|�3��$K�����n��;��[��z�`"9��HΌ�=7�5������w~w!�b>��?{����xg5��l��S��x�B��L��}��791M��.�7��B�Æ�C�Oθ\�E�i�	X�j(Rg2X�d�ل��1�W�R8�!t0��KP.r࿧N������M��BA��\�To�������Ĳ���^4fUE @
�3eF���'�'�����9_(X�S��q�̂4j�q��D��)�(9�
n4f��(HQ�Ǎ�	.5�jh�b�ķ���<I6�����o��A���ط�%VOL�Sq�eW�X�x��[o���xLx%x]ؙe�)yņ�>#�a[[Ǉ?|��Gt��c�s�+�$ŵk/�%����g��=�����L�J��a7�X��X�R���>v�Cs���z_���4{��5}����󫮺��w}VݻwoS+���?z��?���wu�y��A�o!��ٵ�g�~�����V��t����>̚?H��#�������n�!������3��fH���mذ����L�NL�:�ūV��h}c��|vī#�gw4�NSx�� ��2p�����J ��^���%�_��'Ԁ`𤑏���b��/^������+��!��y�M�|顇:|�HSS7Y�������(MG�f2�`q�8LX��'ml��֧>��m���ݍ�������d�,l9���򫳌f�h�U18�$�j��'����1�-bb���s�( ��(0216�V��6�@I
[ZŤGP�uH7�'��44����X��t�a�^�}�C��[�71bp�x|5�h�@�dK�8"/��Ji�x�����p�
���2���U�G��ߥ��!	�D�*���Q<��+��N`�%�:nh ����y8��7Dbdh�2]�F�k<>?�L�Z�-�*����g��x�B�Q99I<�U�O���.߄0ز+˗/����϶����%�*����[�=�����&�e�0XSʃ²9����?�ȼ�2����k��� �u�j��I,�UM�����ηp�b�n)T,vl���i���)����!�
��傣��O���~���ꫯ޸q#1 �%oűq�V�>����Q�{�̰��vq��W�s�n�!��]L>����.Ed<U��[��jIw�E����|m�ӚN�`v�jq��M)�H�������y=���_��ӟ��؉��Z�e�j�U�Ff|2S#VR��N���?u�͗9�w���@�KmU���K�ϔ�e��?4|����;��*�sO�����Q/�7$�AX��+�qlp�8�g��;ϱ�5<�q�.�&Q�PA���h43M/��S߷���d���2ܹ��s���{�}{��:x8%a���
ʥ�����X"��n�F��b�hm���z�)�N�uN�<8��-Z������/�8L�ok7�����Hɡ*q� �L�������Ӿ�ۯݲ��_���\����s��P��R�\�H2P(��b"�Px�g.;�2?��D1����>��LU%#TSnR�C\L3efQMc�\#������m����i8��c%���;���Mn�/MM��"��eBф�bixx{OD�n�?������F�O�k���(Tü�80x4�@�:��%��u�����N\a�u\�c��@�fT�`pYq��i_rp��W���C���Mu��U��tM7-.�ҥ��?^τ]8<e �b)���7k6�9\.U�u��YM���+W��a_���NVH1D�CE	���S���ۋ3�1w.6ʄ]�=)(&�y�zF�,Y��Kb)�uAX",����. ��s��KR5����5�]Qu��E�����giEGm;��k!T"ժ)�81o��6���Kp8 Sq��	���?a�v������Qы�<j�]���gŢԼ�QȾ}��q�#�l��!Q�5�����\8��ؓ��%S���vW
��ʨw�PE�Ë�!�����K34L�8��p�A+�ٳgæK�,���nH^�m_�v->��������] l��ԧ�D�;��n?��/u��]��_�
�
�Md��$�XK�_��3⚸I	�$\����w�T��Y���r���C�Ѳp2S�K�TW'���u���b��ٺ�́��$\k(��T���K\�X�4b	�l�|��JŢ4�Df�fy�9��67�7Q� �vK�'��P\�<bG�k-��He��h�����'Y�r� K��/��r
����t���]!���ݴi�#�~�ր���Py0~�R���t"q�h>�"ʹ�fR��@v���]��s��-Yt��&�	���ȯ.]'QI۲���������m�֭���jSs�_��.N��ÿ�1�B�"l�f���S52n ��5kƬ��~��Rp �+�+�6��*YBͪ�)���ho����\$����K/�=�W�W�&ۢ4d#F�>b��U�X2+G�N�hSS3����Jx��W^�H��G��9w�'�K.�Ǐ����d?�'ۂ��/]��2z��Aآ��0�%���~�p8�S\k��4�����^+74�557tww�Baxv># C7��b��g�}z��5��;v��l�C�H%�k�?y�� Ÿ���c�`!�*Gx|<�;���R�ɡ
w9s�+�9N<�̣�vv�|�����o>v�})���HL���X"�M��� kC�P����Lc�C�nJ'S4�M�1������~��ڱ\}��L(�tC���7Y(�J�0̧?��:Y��i E}{����
Tw/K:K�t f�@eo����4U��^y�*�����C;v
�q�M7}���є&�	� \�Z��:�م?]�mۚ5k����1-joo���o���ry�2,�@�cb�P0���[��=�����@���0���V��tr��eN�p�@�m8*)
R^�(n��(�f�*����RYy��f�f�,�(�
���,⹭�q�p��֭�|�m�߈��W��f|�c�)7�4PjP}����[B^X8�:)u�!��Z&��U���k1m�m�.[Z��_@�����{��^6�����}���d����}����eed���?��?|���UyliE��?(�ү����B-a�$�I�
\��o��^��#\2Ӆ26s*K���.�AK?rO
��'ō0V��x3|Q��;���O��߈g��ҁ2���F����5cA ���K8�V�~{כ8���w߃>�{�n�;�����s)�w-^�X�'�sH%)�'�r��pC�d�b�|ox��H\I�2�*�rŵ�+��C�J�q���L�x��,YV�/&Ր�I��Ԝy��6s��5�U��ux��޽�Է!<�&=��~K��R2}}p��ϧ9"�� ۀ�"��aİQ\99£�<,��}�`��̙/LT����ڵ����cF3�e�D�@0�MM��Sh.<�B���pF͐P��;�}r��|�� �1	MfV�zy�c�x"i\�ͣ��t�M��Gy�߾���F�����W�����09��aap�j$jwnjn��	���i�]&�hL��l&95T/��y�b�����|��|VR�x�\q,����҉+��"�{4G����8���p�zp`�ĉ���R,ۼy3W�9���dE�.�����E!Aq�����&Ӂ�ݝ��m���?��Zr����4���/ ����t��:	K2�-A��A���u_�\*�ZgP�T0ܺm�L���g��o�ticKK����B>�P��o|��C1A�n��V��;{��|�J/����H	�@���}���Ea_���}���u�Œ���+���xcצM[�USU��%6��kO� Q��g����2�����GE��D���JQMw��P��<��i�M�6"�\Vj@s��u�c�BIx�Շ+	O�	��x4��45G�<�Y(�����u���bf	�b��$�\�t�ģI/�MMt6�2�<ϬV�>����gPGhܥ�]/�|�2������/`B��6�D:J��"�[u<��9���G��X���2�lc�,n����G��B�I;�p���<w���.������@L㇉,�&C@?q3z��g��|�r�=�Q>����zӍ�����vL'OHS/4xCc㫯�z���%����Jh�#`����ʥ+�/$eM��U�_=�u��{7�߰q�J�Q �`$"u8+8�6n�tMJ�-Y0B��Ҍ3�?@�D#���֭�<s��?�1��K���QW���X������ɬ,�h���o>�#`N1�OP���T�j���2����yk��_��3��i���h�T�|��;
M(���`!c�b	��0��B�.X� ��m&���;� 0t̛��_>��Ͻ���(^����K�@��ċK&��`KaB�k;H�$4.�;PnSc��w��6l���{�;~�<��عs'v�����
�)�_h����?eԉE�讈�8W2<8@ν�R�1O!t
B��ɡ>I�z�y�M�S���mHL�Db,[��\7�ˎᝀ�R&�S���Ͱrx�S�N�?�#�W�l_s�5~/�F�r����_��M�)�p��e���\]����\�P")m����O:�ƷgOcǓ�BQ]��<����T\_Ay�DXpJ"� n��h/v��˖-��"�D<!���sf���]M�Q+0�P����w��݁�����[�?~�e���|��=��_��W?z�G��7h2�Ӄ۶mk��L���r�X�b�[,�V4�J�i��������La��?�W�y����իW�6E�Je�y]�t�o����ruɢ��Yq��n��G����>��|�՗v�:؉g�y��W^����7����?�ф'���c�\%3ً���Gv���' �|��5+ϼ_���3���ҹL�WL/�l���P$ñ�R��OB�j&Q�&5���p��득�g��(����e�Y�g��B/��Q��0<4�7F�����A��J��t�@�J����.d�L*���4w��yx.?�KH�=_��_�xB(��R� ]ظ2�����K`�N��ul��h�#����������S?���� C/q
�PJ�")�eؖk��*���"�UM���f-��bɔk9���b>�df((�]o�JUS�`:�����>��p7Է�9�Y)[�d�csE�'1|)�pa���C�?�By�I��[���JT!|��&i��C�>�(�n6OQ7�ٌ6]���.�2=��I#�#�b��<<H{$@�K]*(���z�u悎�D����j^��5dz�N�:���!��w�_�bn]�q�\6DR.,``Z�����Q����~��*���3��*���G>��;��������t#�(�hH$c��˗/�n�V Yhi��t�Q��k�\�dZ�����{���H����y�ׯ�v�!X����� �{｟���6m�W��B�0����e)�t�P��'m��������_��K_���{{��~�e�$����!(�R�%޶��
�W�V����<��n��6�)�a8���6��9�Մ1�5�����Xi���O�_�����[nn�Ғ"�K���1�ӟ�$0\3( �5F�,�
%������?� K`쫮�J�=�n�;���ˑ��oߎ��u�(B��g��-��s�0#�c�)���I��S?ɺOC�u���
� ���fb脡D���$��RyB0e�bԀ3ʖGjs��+@)���7�ф�KFۅ�;�)�Z,b��x�P��+Wi6q�J�uʠ�DA#��1��3g:�����R�Iŉ5j�5xI5�:K�������LKI��M�L-��Eq�vMO�-iX�����Fh��K���U�)8�CL���n������jYl 8��0�P�>�b_�ĉ(�m�]��;8*w��7X��|����œ�f�jCM��[�:�}���^�f����>�
9�ƈ�7�i�Oq���?�cs��و{Ù!~7��t2g)�%ׇ���o̝5�d/Lѹ�I�����1>66w�\j��>V!M��Ҵ��7���/@��Ξ=����w�ml�����?�!�1�� '^/����b=��_����Z�H��̜Ur\舨V緵����n�4��V��;�։Ie��49�xr��2�ŲeKZZ��!�Df<����?<6>~�������w�uW{{;�]{��Y������T*�������^���F�(����>s�^����^�v�[� :��7����J���F�?|����_�~=,'�z�C� .���Їn r������w+5��0t��J5tW�v1J�p���"C�;��
@��Fb)�a"��;�k� ���(t��x�����4Q �J���U�766��Q0lh�b|4ƍC�/�S��ϝӑ�r�L)���0�PƜZ
(�Yjlj�
�t���+���F�An.��9p	ꗩ�oNs��}fT�X&��¯*V�R	Hܻ*��P����=�R5)�x�����f���W]��(��@���Ε�4����q���${�ޖ�	O��}f�2jX�L�@D��s�3��X��l�����If��o���D����/[���ĉ����P0)�}(���f�: �t*�Kc�H��c�o��4�p�pw&�BeP��۰�T;�s�/�X�TM�����>�Z��o<�{�Z��Ʀ��k�(.�WY5S�MS���H�� ��O?�4=���\�K$p��q�q���q�����?�w��p:q.�"����F���4DW��fr3[��?y࢔S
��X*a��/y�"9x�{��1X�E/ټy�E�����G~׮]8[�l�#C����\g'$��K�=|\
&�9�k�
���?o�T|� ~x�>�<>NdO5Cb>�{���q)��J8���)]O�Up�RQ�*;-�M��X�����F�`�'�N�(��g:]�g��EdXN6�Tj�֩�#&&(�.366m�(�,��������{<�_���94\m˖Mxe�외`WW޳j%�rP5
��7������E��Júr��<�\��C�A��e*v�R���G����[�W���z���Ɩ �?>�{�L�N&6FGk�,��[?}	����a�U�*N;�WI%�D�e�ԗ0	�j��>zr/>�C"ч'NbB���9��'M�0��������{��ZF�>B���L7���$���D��g��d����Z�jq<?1�i���sx#����2T�A��d&N)��(A��9��Xn4��7�h���Ww�1>2��omIqcv��5��?�,��f�b��'*�Q��T2IY5�jn�E���5&��+/i�v�m}�_��:\�:�c}V1��/e�������=T���%�FF�``\x[GϜ"��*�NS)��#�_����O?�'��������^�
bD�[��_��Ǧf���ܹ暪��;u���#g��8s�̅����в��ރ=hI����r$ ��a&h�^����}f��8M[�t!�1�y�����8��LBݡh��NOl�j$���y�8'��h�
�ǃ5׉œFj��XL5��|���<�r�}E�����T������9��X~��)���\)��2#���UO�j�:46Z6m�:��)�|}�+F����ԩ�+���L,_�\X�<E�Tk{���=o��l�j@�8$���n�)�/��Q%8��� �SrT��d��b���� Ք�F��n���]�
E]��2y���j��={��v_O����~���[���:0�����7�t���{�k_��/~���9��U�J�H ��
Yï�r�%W�.Ж�ё�<�Gj��:�������=c#������w�
��:�f8���!�J([,�ݻ���"�sY鈁�!J��px������B�4|a��teҩ��F��LS��$� AU��ؘ�	�œ�\�酞�fTh<�]#5�YB~W�RO}Q�gT91�*%w��MƳ����D��'��W�bW6Q�ҟ�����nք�
�L��\Ĉ+PB�Y�T�q(,_���-�aL�����hk� �$����x��fЙ5GjtX��$�@v�	`��9-f�B��ۀJs��y̩ɵ*O��k*<7��g���G-K�#}�R\/&��o���J��tg�(U���R�*�XWq��N)@|���N��8*J�U*yKL�(ġ"@C�C����ɢ�,�7���%)8
B�h�M*�-�MxFS�2Md*�%Ә�t�gK�ƳEh.b0���B�sJy�4U�x0��dC)ur�Ж�T��yz�n�a��7��Q4���il֏�����Ǔ�.����9�%�P�`SAi�HL5'�q�J�! A�各� }a�M	�(_j]`>����yG�ř��P~.C�X��Gi2��h�d�[hjC��������*�z�3P��08�e�	���<M��0��`F�IX��M�(U��&��&�	����������y�.x��uK��~�p�����@��� ����X<t�Bev�L�/���Darr��Je��!�Y���ؔ�|7A�P0�J�|T;^���Т
hʭ�3x��M2�D�4T�φ���L�h��K��j�p$ʵ��G;� �˿p�J�@Xq�ͯrQ�!�n�d�(<13�8҇!�G�LH���F҉$6N����J�h0�}	Pw~C�`�B�X(HC0�;::��J�]��|�0��0�v�4WU|Պ�D���1o��\56�C&��1�#^�L���;v�pq���M���~FLq�X�r�R��¼���JN�cO�J����r���]���#7�gJ�T0�Y��@b19T:��4���y�I^����M���k���7���М�jzނ����O����+.[�j���'O��{>*���<��c&(��QxD;T��X"*%�Be}]��n�#~.�'}Ua�$�F0H��,��T�b�
*��ts�L�T.���6��-��N�)S$�Bt3|�C��W���9S��*� �_�(�g:<7B�,~�'�FD$�R�R� &������B~PJI��u�]�1>ָ}F����p-����:u����H �Zf�Jc�D����CS-R�lZ�k�|lbA*+K�ȇ61����t�����ja١�D.
���=!V0�*�	�I#Q�7�m&J�B��y���	3U���NֵR�,�5�����,.j)Kj[0����Z��-���Ir*=(����i�2��$��g���8
22
���:ԩ�JlΕ��+a��ċxF[�����\�4|1��gϞ�'��v�&��ӧO�I�?E_L�IrjpKG�i�I� �"W��2>��ɓM3Z(<k��ZR�H6W`zN����=ӊC�̙K/�4R׈S����FUT�V\�v�]��,Y���L�a7{r�pKܿ?@j�a�$˕Z.�"�l�-��E)c�0�:e�l��X~�����7�3�@$��2C.f���z��HȆ�δ�U�%2�.$̥r*
�xw�߬���_��u���dja�U]	���
�>Y�D"�ee �P�K�$�8�dܕ�RS,��ߞ�G�m�ٶl�F
�ܛ��[�pn"��Rܟ��u;#�1� �'��Ґe�dК��jJF�(�a�)d�i5�R]���ZN�R�W
ĩxr<�����#�l�(1�%Cq�H���`��m���/�O7֑�P$S�)���&���K��f�_��*��! 6~�+�fs����sf��3�/c7aZc��.���#��Ц��b8���M��aZ�8���3�V�H��cG���2��
���|���Z'�HV�%Jp�R��\��!�$�/���+4z�jf���pz.��K��Z�� (�AlǠ	4�k�jT���j��ժ��]�)�R�Ui�� �xX�h��T��W�D[Qa��W���5��[gu0���\�xG�疮�ml�hi���Vb�8��RW��i 
qbi������P���ġ�s�Vk����0�'�9j���TJ���H+�b��r<_.W]�|���p_���Eu�H<���@J	���i�� E!�&��3��Luݚ(`���(� �v��>m:����2T���`&S�{T����I�>P���FH��w߭����g�zM8�_}��y3n�QB>-�$C���:=!u�x%���~�!c�Zx�!r���+�:�����5��/$�b�'s��RUJ8���dU�!D.�H5!zT�A�Z��1Yq����b�h�'G}�Ib�NE��ȧM���N� [����Y[kjT�Whz�iZ'��8[���p��Od�bry�1��656�ݖR��:9�K
s��Պf>|��2��X��T���Q-�e�p�\����1���-4w�,�G�@Cb����8�eS�걧�f��lZ~Z:�a��p��M�n�L�ѽ]��3����	�'� jr��X�t�b��J�j�9��g.���d�`%�y�6���J䘙�ƃñ�7O���J��!�!�P�U����#E6��R��4n�Eb���h��%�ω,1.�~�t(��L�񁱱Q���[@UTqgST#��1�6�ׂs ��P������qh#`�����Nr`�j,�/��5�R��2�0'�[�l��SH̦����>i��g�C��B��gSd�sU�0�EC�;R�:Q1
�:<���m�JN�+q�V�^k{;%� j�u����X4D��d`N�����@�.E�=����uJc���AorFwU���6B.
�SJ�iP*/W��_�ߚI��+��OW��7��]W�z�~�a�hA�L$$�V�x�Z� Уfŀ4|M͍��8ސj�'"�=��2I���ŋ�\��(3�I�x�*?nh�pE(h�}Y"1�Ųk��"���W�p�KpX��̏%S�= o#��T@�i)�_�i!n{���?���7�5�:q�����-msLG2�f�B>
(P�~�R�HrL�Z�0�rY��]#��zUX���Ҥ��x��h�8�����`i��	��|A��"�N����(4��:���BI�U��D<�e�UU�^
O|Bu�fFf�ze���l��62�n]u(��Ӿ��Tvi�<��2�s�XU���u45�)Z-��jn����%0<
����
��744�}�v2�TקJ��|	���^���N�R��Scn���Z�(��du5f����0�b�wa�f}I��/�3��ig��\kk+<|�b��+����Ķq���.�h�"��eUx�Հ���W�/^�7�tq�m�ƅ�\1q"�S����b3�m�E��}S4�E��󁞫�|eC�����t�ر�G��g��G-~*M5+��;�J�B)b����BT���,B��w�+?4B�{�"�"rIou���]�=���Z4��[�w^~��\�[�&d�8H}�X1J���e���\*ɏ������IO[��p5��spX)W�I'Ԕ����[�&�\��� LFV��w:� �{�t��rp�aH�4��3���T�2��E^7��,>~`Np�D���2bg��H��b�56���$>N��"H<C�IG��#}�@�����BO���u$�.Dt>ݰ����"��%B���jl�K�:�&}�H��i�}B1��P8O���x�����	G��k[�-�L��lvB�p4T.C�A8N����h4688�E�Hŷhђ�P7~���\AW���Ib0�:�O��"j>cd���8a�v��~ϙ5��K.i�;��ɓ8��|QV/bw���q�,����a�N��LB�::�͟?�:���;��d<v�����hV�N%`�L`�)�A���s�fT�ܸ$�l���ST����[7��tO�W5-H5�-�<p�r����W}p+M��R�1�2��n}\<iڞ���;vM#j]����=	ZvE�a1J��g��XC�x&�l1�p)nL4]4L	k<2`'ԟU���DAl�|+�@8w��k�*Ώ
����0�X�j�2�Bq������x"�i ��E%t���ߊ��j�A(]���?���U��}��__*���+FF��]	���z�g��(NU�:4��rB�\G?��[/��Zr�����Lw���ߏ�"���B� �&�� 1 ):�8R�!
P�gj��G��|��v���D������8X2�Z� �#4��L�l	�GQ��ckq� ��!�%z.���"���b�^����G���6MV��ai������Ťҟ�U�z� �>����}�c&���ěf���w"�Y���@��RXM�SO������~����p�Y^h<����_�u��}]]�͛7�x˭
�֫�fw@�}�Y��Ӷm��B%ǀ��sA@ ���ꅋ���lC�v��ơ��oji�U*�C�1;}�С|vB��L��D�ȈCα�LN�c� U������ɏ*�o��S��~����Ä��8xC�.i�c����Á�ӨIb�H۽{7��nL�0�%H�1|��������_�u���˅z'��	��V�Z��(��S�����#'�������+�u[�lY8BF�R�`��Fc��Ο�W��z��y� y0~iƵ�ɘ<Atͨ�U�zQa��)_�T�&+V�x뭷�v����F5q���	��Ǌ�J�D(�grձ��O~�c?��ϔp$�r��������v�x��],J,����W�9԰^�IE�a6G��3��9��CE�3�zʯ�J4^�1n#	Ԇ8�Jͬ�.f���oKS#̗��-�#�����`��ds�b!ǚ8�J��j�����szw*aF�MǙ`I�yh��l��JGG8�,��|��?��f����\7�����3�I,��z���U�{�N��0%?��+W�:z�����w�z?���k�}��![��
;��O�l}�3��.��������/�r���K!K�LN�q��JK��uu7���b�b�F�wgμ���.�+��b�ʕ8�8pX�7^{�����o�q���:;;��q'�|A����*��N�mk<�H�\�T*N;�"���o2��W/q2��>�G¨���O��|4F�^�fє�j�aɨ,�s��2N5�蓸���� �-M�2W���0�y�3�<Fv5J�6�jٛ5k�{�9��F��Ќ�`4
?�R�*<�0�d���8t�V���y�kV���'�ʮY�B��i�?kղ�$ oيC#oi�<.8J����Ym��͵b��ك���������G�-�i���C@.k�YW�IN�������z�w�7t��'���\g�p��ܾm���O?�4|�x,���Q�AȶLa��Z�@Wj��:����B�hh�֭R�Eó�@&0s[GS�Du���
� F�e�B(	8�4�`|��U�yZz�r`��*����I_�V�馛ps�?���^�\�!�BϚ5zBr���!�tlO���mlL�w�}�֭6�Vṡm���f<#�dɒ�)^��o;�7�ѡF�(���L�=�����8dl͚5���ԉ�a� ��_�ΝS� x��{�ɧ��E���t_�9H�h1w���1,�T� w�p&�<M_�/*��/��2�gZ��E[a����ٳg�'������$=#	X�q��KSu	����B@��2A���(yN�B�&�0J`��<�9<��O!ɒ"�"��G�l��#4��$ H��� ��Jb����_�)H�3�ƅ@����ai��x�G�m��1��������H�ƕU��.�'�X�[	��Ã�2%"���a�ų��f��o,̫v�@�a}��uA`]gFۉ@�T�i�$3D|�r�tr>�d����}�ݸ��ۿ}���y�w�1w��o����# -�����[Z��P5�)�gV� -3���?�Ⱦ}�r�p*� �
nh� �7�t���aaǫol\�z-�u����t�K/�t���8�s��ڿ��Lx�M1�p��7{Ν��;V,_���D8��.X4o޼���tKk��/���s�}����3�"�8A�x�(h�D�w��y��~��W��F������ToeF��ݗ
6p�#����)%�Ds�$�?]W IR)�������A�uz���%=1>��c��%�Wn� ������[;�ΦQj�μw��tC����8>:8��d�j�+����?�k>������K7K ;W�Ԝ�"�x�f��ݏ}�Bqg���_�"����ݽ�Sފ�[�r5�B��C�����"q��B� �/�	9m�(�|�H��܈ K�����1��f	0�Go�h�G�	O1�����E(N]���ҌR�P^7���gq��P�P�U�Oap�4õ���om�.
I �v��0�v��'�������_�4�>c����Ȩi;���p�r�Z�ա���Μ=o�B��s�/���.W,��s�ը��/}�S���@�6��!�];��x���ݎ���}����W�����y|2'�(������d�9�G�i���,������C�E ��B��_���=:�ޞ*Z���R�����+��l�uScCcc4���g������o��l�C=����g���5�9(�TYG�<0����Ϲd�2��cG����$�C ����6(��{��~�i�\�$�0�@Rjp��	�V�k���qx\O=�,�fw����?���~�j�"���~vccz$Ӎ�BE�n���Б�W�S��F�(;J		"j4$R���ڎL��Z���]4�T�	5zg�	��v�\��]�c��g�6��i�Q0�x�h]��I�f�C�K��jƗ~�ӟn׶/�&�F��$�d�5��_�?t�7܀����C�����S!�\�=�Dw��GL��@����צf'�\�N1P���>D��-'��(Fͅ�k��'uj5�0��1}�:��?�
��g�� Rh�ۃY��M |���GQPM��_����	�4G�������r)��|`���F� �~�5Ǉ��D0��K���dn��*W�a^����R8J����  ��/3�rRo� ^���\Zgf�䘑,�_q�m���*G�]�S1:>B�k���|�t���5�\�z�:|��'�&|�5Y�x!��7��'?�I<� �m���F�U4�-W��� ��.��r��9�Z�<�#Q��CG��.YL4>XbrHT7[�B�[��qdq�������#c�n��=�p����pSc3�,�#e�8�]]������.�͍=��ԅ`N@'u����*��n��C��A\fs=4�x�^�vm���JՕ�.�%Z�+*�1(1,�R$�<���_�"�ZT��-!�	
�i�Ν=��|7���j��I�M��:������PQ�Uۮ�on�d� �ͭ�X���=���~���?�<�ڰa$0�H>�ԓp3p�t2�U
!J�X6wT�$	$�L\�UpCᔾ+O"�2��ٴ�a����c�\]�~?��U�=�dX]��0����T&S�:LL�s�L1k�Y�+� ����d���P}Di��K�C�Z��L�2cRځm%����8UW{���`owO�T�'�>]Om"�/R ��u�9�g(ަ�.�z	}�@�R�� nd �4B���$ʸQ�N��8���QHBՔ�U6��%K:��p��Eǆ���`З��T����K�H�pv�O�U��������T�S"��:��s�'Ɓ�����	|�-�܄��M�6VidhH�����7�Z�b�\I��C#�����=��?R+,TMӃ�Mw9 � �n߾��E,W��?�A�n��]�bţ�>:4�+�^��ʦFJ�n�M7~��=��ҥKq2V�Xq����L�ػw/7����u��_�j���X�����[ �F�pbJn��} '�w��/FF�s�����5}�$נJ(,!f\�$��:?H��6m��y���u����+_޹_}������밮0PP�@�Hx��[�g\Ta���ﯿ�:;{4�b��EЬ��ډ��d���{����ԧ��Rq:?�O�������4�+|RiD94�G������$("QM1�R�/u��t�� ����fIZj����Vף_�\Og!��J��|�i��P���_�`1�4�4[Rm-�+W��{pe��C	٩������v��,0�R�"ay"YX�)N��
�/�d��R�:T�{���!���U�8<$-Ū|RF\d��"�6������Q$n���4<50`�^jD�Q�����ri�����i��P�2��uS{Ja"� 8���wQ8g�r�86�E�Β0� qVe��O���Swft?�Y�� P^sCs{s[﹞h8�0��LD��R�m<~��Q���`3��*��J�g%��V��s����w���{�i��EGO��?�TŲ�?���wv���0Lx�\)�)<���e2�����׿n��������g����)<��'o�zEGǚZ%_��X���S�W)C�G���ZUr����M��Q�P�LA�V����W^�*�	l��Μ<�v����f�u`fH�ʕ�s�-�������70<v�5��g�2��˖��}�]-��g��Y���&��>��#]+�s�[W�ۀ���Wl7���c�d]����m�j[!�}�g��z7n\_)�/��4V���d*�P0�v,�\����|A��A�f	�l4��zq:���ê�A#fh���*fE���x+��R'~���qL��M�b�bt���F51�+V��\�Z%��.\O��n���Q[���P��CC�ga;(H[�Ujd��lq���)J*8V(��̐n8�q����晪[3=�H��N�(�H>�.ݼ�f�J}��GF������Ž�O�K�!B I�v�H����F��uh�J�x�wqo�~*ߏ]9y�߉���B�����0�V��9���̝[���y����{�5����
1�EtZ�\c�W<}�4�8~k�ҕ�)��O�c���z+��-Z8�Z�ZZ.��{�"\�tL�f���7���Ǥ�1�Hը0�<��v�`��c�*��"���p]`_�a������F� Cz������?���l�u����~v�С���W������_}�w�Z�gb�&�)M".f������+�@�C�d�� ���Â�۲Qr��9�\Ľ�&�O��I�m��*'�'�����u���;��0��/=/���=�ܭ�|߲���P���z�UW]�5�x���j��H�������~S��A]#Lg⹰ �O��/�6m$^�Ƹ��]˪d3��H�,΃y\��y�>5؍�'��5�r�Q��gX�j7� �T#)m��B�t�[Kn��ىӬ��PE���ᘹ�XB�#.�0u���YA)���,e�H3cC��,��dq�) ̅{��g�$�;��+���}=@Rs+	<����WIr��	K%SW�ʡ�ϟ���/Y��X�����/�鯿a�Kq{2�
1dc�p�=\*�w�}�p�����i���]�Fh������w�����±���|>�-�W��������{��Ξ�Z�h��S�ƚ���w�s4�8(ܲU�;���4�������r)	7����@�VI֧�.�s��mۮ\�f���cc**��rJ�����|]2��(p�=_���"H4�kW��1̀��K4Z�
���h�\�Ξ:G��N%�R*r馵����^�qi4�s�J.;�X�֖�T]C8������J��j���b	���žޞ��b�Uܺ��mZ�w�b��'<�M�+��iy����!K/�>��s@��T������/\�5����;Dy��q|4�϶���TR�&�?�����#��Hĳ���^�V5ԥ�5�����(D����P��T�x,�2Q�ײ��D�aG��(Cs8=H\�#�4� �B;��	���Q��h�N�L-f4J�)������?OF}0×�khmm����"-�.Y��?������HD�� ˳�4�Ul�sM͠��ișeג)\-E�J�dH!�-b��<�N]74K����k�C8� ss�*Ls��]x�|AZ���1���|�+5�O<d��/֜��%W:3|g�v�ݸn�a�eQ�b�������t=a�K�u�-L_$��l�ǳ�,q���U^�ܹs �=�gK$����IN��:��ÿ���T���i��g2P�mni5��m�Kc�J��<��w *��|�9�
:vOO��j]r�%Bb)c��{cC3_4AJh`` 8G��^�wS�W2�F���F��+ܟ��R)X��b����:İ��3!�'�/�}�hâ��P�B4&���kA2Ԭhi`H<N����3g�T�����#5���gN�:E	��z�pkk�d� ���_[��L��*ێdL&��a,�"�}=��ѩ������h�&1e3 ��d�V&��n�q ��6eF/DH��X�d<�H��O��]nXDήOvNy�y��JgQ���R��0&�'=)%�%�ފ�ߛ��dRXujj�t7�x�pɠ��X�T*�Io�ظ�6���rQ�.f�^,�$cIW �p3�
���G�&K�&�S���e"�DW�.�D��{�?J��B�*t��f_$k�2������@˾��̹ni�����`=X0<�ߟ��2��r�A�y�,������o��?KQ��W_�o}k٢�XX<Λo��ېzI����{�'��7^��[ba�sZܢ�3�{�`�WW�8])���dbt|�����S'�q�8>:�|����B�x���m�n�3߳p��}{��e��>�X��N�=������w>��<���_�򗫕J���_W��]w����~���o�/�&�ɦ�<j�	/J&u����$�tl�S���K�����C���hJ�YC����0�����5�s���mZV�2lе�3[�ŌY-E#����8���T����>�9�)�����~������f��.�T�d�5���`�fa_��V]u̶��z��m���Z.����ɤt�ǥV�<>2*#�p�I��0�Ԏ����ed�������G�U�>Tf:�p��ͦP��o��"'�di��8�"M�4�AB���=�N����6���,����ȑ#��8Ls�vD���e����j�,Bp��=�_^�f���ۙӖ�B0=�g�>&�[4sf�6ڶ-Ӯ���9�I��$f�������
�)5�r��ȘĄE&�:\�_D���^|�uی��Q���a�+���9s��XX�P�R���c��������r��˲��������?P����l�z���{����o<�.�ce
h�VWW4�9�[s��w.�d���][6lnln>w��+���~퍺O)W�b�
s�QxUAܾ!y'Q-x�W^y���3��-�ͅ��������cG���4P�T������!�AB��O|�%F՝�O/Z��F��} ������bk�p�)�c%�������������]Y��b�ic�i䇱��xJ�J	�D�Lu$&x�*�0����|����U�+pjq2�k��[DwB�N�  �L���BX"\[b�t�艽���!����<�`SZ�%;OU��dSj;�5�RT����)���m�*���-g����S�tv��G��6�uR �����:��N��I��6�#���R�*�\��0�JI��C����3��Ʀ�8c(�j�ɺ9'�8����H0$�"��J��|U��K�)� ��1Y��}6b�I�E!��.�}�"�TωA��@�Wee$g�K��/d2��d��m[�ھ�O��?�S�oh���]_��W�Μc�T;����`�"B�Lt"�	O{�G�_�w���e�b���j� �!q��#�+H�S���[W�p��q!�	��c��h���/onndJ����/��"@\R��+��\6�kʉ�g���/\���>~���F�|���ǎ�_������n2=�8y���4���kɌD±�kz���G(\�L��Q���Z~�������Nt����d|�Z)��f�����1��ᤊv��}^1+4�=�n*�4�(F8PJƩ'��"�Tt�O�s�3jk�}&g޴T*���j^"I�l����&v".��$E�B,����%[�<����Ճ��t9��%� ������0R!�F�?�4k�2t��^%NNإ�0���0 ��p�9��I3$�e��¨�$�$_�1�TNJ�.4�����ى5�6̚3`��J#���c�7o�L%��#q�C�r����8p�X@�`�����'�T+$��.4X_� ��m��,��fr�d�D-�8�e�:� �W\q��i(i�J�'Ntvv�8qK��>Cr3d��\R�T�q��eZ����V�=���ރՉ-�#-�8,>ũ������ج%��%%�s����R��e;��~�U��e*X��_��>?�����r��,�g���0{���k6�onoueG�xbo�!D����P��'zzj&�}�\2� p��i�q�3ϟ�p�[ �Q����V �<����yX_��4�-t	��������˄��O|�����馛�Ν+*Pbk��"kJ�Kxİ�x'�Q:�o�����-����Ϋ��g���h��d��Vߨ1%�L��jJ(/J���s/�'�E{F�ҝ��-��RN)��T�HTP��qm�&�p�d��,�N,���9͝!�VU�9N-��hZ�C�����~�#%����۷e�t��$���L�nP�)"Cj��3��A����=�9!0A��Y�9�1d�,�j�'����P¶�}2�Jh8�G�̙3g�S#��:S���^w�u��%�sTM���ō7RA��Q��_�
i�/QKK�� G>�5Ƴ$NCQS��q��ĵ�%�b�%�*u���bD,�� V�@N"�Ÿ�Qf=;p�Z�g4-g*^���x��앩X�a��N���ѣWn\!��X�K7^
���w�|�O~�GJ�ҡC��g�\�b�W#2�LPe��0.�E�1Cc.��}'9��zҀ�sɝ�`	#� �	�o���.�noo��GN��niiQy�@fl�_����_g�^�w\��݈E�|�r���L\}�6,��yv��慞qf����8}�4�$w�m�X/^>ǣv.��.�Ι;{��0�m��ݻv�������EG��VKcc>S�CQ��3
QQ��&���\!�b���2�/��2ϑ�ۼ�)����wQх�V9S��xl��ң�޿�i�ag�+��zP��-M*�8�KI<���REe$&B��"����D߱�F�a6��%����"��<�k�RLf��9X�����
��Z�|�؝r��t.<q��
\cJ�t�b.OC��A��J�����]c��b�H�;$kT�j�Ѯ�����H��	}�K����a.���gd
�����92��o d�Ho��|AOm�X5i:�pL����+�e�}�
�����5�[�:wv<R����I�<��U+Ǐ�[W�M�Au~�����1E�˵|!��M�df��o��/����ϟ��ݎ/z��I�G�V.��C����aOaq�'N�Z�xi(���r=��z�M�P(�]�=�T����b�����|��(����<<7T�X�s�=�`����#z�|��ݻ���_�#�oq�;�U$b�<m���T��nݺ����m��6wn���4���V
�=��g��NH�GY,���2���nb�����v������
�p����x����<�W ������?'��*�H�&ӧ�Wi9�c-�>�/�Z�K\^Ψ�^��Uժ)11��g��zR�!��͐�Ir�s��Q�p
W���/P�ʙ�ă\VB�VurQq�lL��R|�� ��`*����%r��S��WM��p��7�v)}�+�
�+ڜ`��p1����#�	G���R&9�<�Yd&��UO���8 �L,�d��ZXjgӧ�-��M���ۓ��D򅚕�KQ4A'��@,{{{w��a�����dT��;��q^\$��
ǟ�=8��L���J̀��Q�A��ul����;�氮�{`׮]0�x3�bww�ɓ'�]�,��Zx��,e@�|�&����+��_!YR�Ilk�ǼP13�Xx�gU�Z�z����Tɉ�z��c8ʆ"��4
O3<8p8��J%�J�����#<�i���V����@�篆�8uꝱ��4�����-�h���$|,o(��=ڻw�	j���%���3g���;�R4ʔ��W�1��Э:<-�S-U��nqN��5p��*U���R&���,Y����d
OPI"�\�.��Q��~*%����@�*�>#$ �Ur� -�O��4h�H��r�> xB_6)Z:�<�%��+��d~=e� �c[�e ��&���C.��M��j�8)O������89:,{�����(8�{��᭦�N�)'V*V�z=��w��S�L`a�.I��E�q��w�	�ĿR�qJ�R�G�e�2�2�]}��7dmqQ�l	�= ���R�c���x|b1O*���sY+x5��X�xOG#[�]�o߾��!+`�r฻��Ĝ���o�w>��!WM:��Im��/��8�a��V�a�t��G����WnY�я|�Wv�u�]?����)�*�Y��|��g�/_�G(������.�l���N[kk���DX���Ν���s �˖�ԍ�xF������4�BWL��E�q�RCԑ��S�U��d�`Br�9��2D\�ӟ�t���B�}����'���̞M!D�)��K�<&�F�Ѐ��
�ԍGhF/�8a9��[,�⎔JՑq%�V�����Ͼ�ߋ�@�I��B���p��8)�L�<�9s��K-�H�MG�������/*��d4��%����&�\J��VH�� >!>X,�%�+!M��VE�R�g(��p��N{�0)��+��5�P� GY<	�a�6�v!C�+�������9���/�LQD�@��PJ���n+&Ac||p(H�w*.�֛�<4� ��V�ƆKc�j�YU�� fQnى'}ء�K;�X2A�`��y�)(�J]�8�JT0�;
�qu�����g�4X�#��,�8U�`vezC}��2��<�8��Z�j��Ϟ=v���4�C=��/Y��C�?���}�+� VD"DTK���������Ԗ.�!I��D�U`Q����?h����v���� ��n�b��Hh*	Mg�Y�g�ģ�'~�X<R5�$�V�:1�ת��؝��Ñ�h8�.�2;�Hc��2ZZ�*%�I�:�!;��6�t����q�B�p�2;;ǀ�e����[6�{��} ?�����k;^<OeV�iƬ��K�Q�P�Gpnǋ��`���BK���2���Q�K�d:#�9��FH�IH!0�m��/4I��X��q� Z�P��O�#�|�R�7��� IM��W`�&���Su�"�z�����K�����Jx�<"�BN�)YN�d��T�Jۈ��9=��?e@�>��.��t!��B����G�%���	��� :>��dv���&S5k���z�
)h\�+`�����bW�E�?��k�t�c�]�OՅ���֓sH�8�j�.%�/|W}}#y}�+^Rf��~��C�F4l��-Zv(H|�ʵ�������xa4���m�԰��Q�����n��.p�^��٤8*�q��D��?��O�Ν���o۶��9��L&;oނ,�P�AUΜ<���?:8�y���/�Og���R�>��BߠEURF(���Jl]ԉ�愫K�7�Q�ޏBɑ@h��v�KZ%΁Յ�E�4x����Y0�R!n�')��j�x,��?D�˳��؋�,���u��g4&^~�e|��7��Y�/���`4����\3@<\�+��BF؋�6�@__�#�D�Z�*\2i�t��Q�&Gu������t��4�%"G��c����f�G��w��ןw16��q� L�I ��H���ܹ���+}�W���3z����'��=������!�<OK�6^�G���ٮv���D9lB���,u��-eƶ��!~���)"�����,<D$ۢҷ�z����w��Ѣ#�ٖ(��@�mP��
HcLx@ŽD��,<;[�f�O��Cع� ���.}A|"�*�B��BA>�����I}�F>���y�����W<�x��0����X�,q�5,"�b�������f���<��GQ�9������:��+E�1�H��`t��T8���5�b���G,^����n2�,�u0;00�K�
��T�g6�����g��L�"C��w�������}�1�YР+V��R{��G�G���x(n��q���B�b@Ĵ �]OO�U���s�HE���v	�K"�	�QavY�|�aG��r���Zc;;v���נ�]�	GCإR�B�4��D�A��n�Y�	�S*ZC��s���P0��5���o~���k���Vv�,����}�+������J����·����jl"���!=��Ќ�8�����>�g�@ p	�|u�x��0@���V��.�H�FR2�Db,7@rآ��V��Du��UX�C hvv�B,	P79�.�#�*Wd�f���ͦ�H{Qd�9��)�%���:L1��Y�.c	z:�.�?�9�
KB`Ӹr�Y�G�-��|��jr.��h$��H^��C�0fQ[U)���,��#J���4�u�ҫ��78��c ǠFOW�eY��O���/_�F!"ď���0� Vl+�R��.	���Ȏ%q��9��:�a*ǑB����:7��"�x��O�%�I�S�#���Q��J������J�/�`���\B����]�v���_�e[m_�}{5^�B2� .������������Kﾽg׮�h���wuw�k_�\�?�Q�TJ.[Ɔd�{B�����͙���2�Tf�*��M�M�L�)n	�(K��%W�X.��,8�G>ԃ�g�3�Q;��4ϣ��Y�j�9��N`LP����ȫ�$�I�Q��nF:g�K�a&���W^y�Za#�x��6���W]�g�|��-7��{p'�I�R�,23b!lm&"�r���ͮ5�*�HAcի�?���DY��H"�1����l� �UjU�L���x�S�|��u��l&�Jf��W�o�R��ăa��-�ien��b��f��h��e)k,�䊌��I���Cr�XV�Q�������f q��F)�	��UFC�P8��9��$��i6j�E��-m1RT��
��N*��e�)/��¸Ԥfy�	ڪT��JϣP�|�%��-��
S|〗،���z�,>�-P�I,l���3#4r��+U#�$�0>>>=]bV�844t�u�5/�p.��띂*,P�xҟ�����e���cO�Ԏ��P�n�{���Z?���#�ɖl8�H=��Ǐ�[��;����s6���a�x흧����g*��+�t����Hd�<��X�Lɨ�Ѕ|�G��ݨ4�AKy�b�飶E���O^4e(7�q$SLXсb�;J	��i�mWFC�����6=7Sw2қ�b���؅b~Χǣ�Αa�PN��F�$�_����L�P9p��?G�.}�d4��C�y�?_p�G ���<��{Rְ����I�P�Eqɵb�^*�u�H b�]�ĉ�io�2O+(q<�):�Ǫmj�͔<lU���@8��ؒ��n���Z�*W83�����؉�D�[U���	da�`�O��v��~��,��k'�:�"�ht�`u�r��?��+�V,Ruɠ�n�v���TPm��>5����Zo�<+P���9�8�:kᓖs��H�[��FQqI7L��x2q�6�=��*>�9�����
U��H�����R��'	�p�"����p�j]@\H�HC ��jb�%�$�;����S	��43�Qo�ϣ����
yj4�{(��W�\���B<���R$�wǧ�p��\�9�O�L-�g,��y��'�%�ӰQx^�������P\r�lar��S׵J�U_�3:1Q��Woe�����׬Z��B,��O��>��xT��j���rRCT Q��d��2+&E�7R3��֪{��+؅��A� ڪCVM�Y��Rẜ:fp-W�wB��Y\��+P*�<��©SHc�k����O�A)�� �w،r�U���z�5��+
�
g��k׮��TGG��݃ǎ���yƚ�m��t�������e��{w���>�s灿��/-�-{��%���P->ȉ��J �>�{��*�AWu��"#�)�Y�3uМC�b�'�DU$VFs�w���1>lf�|
9~J�b]F�J	7��IgU;R�q2�Hۡ�Og����I���%�ak�(�5�8�X�'�c�D�M���^���)�m�lh�Q��YddBN���(�$��Tש�q��	56č��� �6�I�f\��W'���p�D�G)rqD�纹�D�Ac|,�\Q>H?�YHIԘ�UeU
:9��BH��?F��hEf-D���)	e�dɺ���_��>�ikk�����b8 ?��O���]�ݖ�ڰ��p�!���B�)>�e��$2�NI��*rKK���������z{{Tr��9v�бh�	'S����#�?���<���� ͬ�it�*�"���s�T�=F1���
�9��p.��c5�����5����a�쀳�@�3�k�.HqXy�,��A�=������k�"��ś��Z[[���Ӷ|,�IK�M�(�B��5|��+�}��S*w��Q�����u��5�V�!�������/;3�u���7��$�ԩS��t���T��D�h�B��!��S��!G4^��U�+Uj;�u���W�WL��X��/0}��YTµ��SB�#����q�D��>Idl|�[3�EP��/��c�M���L���Fj�FGA��E�#Xކ+�D���v�e�eJ��Ju4�>���0���Od�f�A�u�Q�$�c	}�H�`�)Aw�RJb�y7d�l��<�j�f� ��c�Q�����Rj@qé��Dz��g�N&����7S�!�t��8��8lF���t3�_Qi[w\�	n=��UJ�PLZ����T7
Tw���V`�5W߱���Ƀ���˅�~��dZ8��XE��pL��lw�������|��5hz�@*��@��zYY.Ҵ�ޞ����Ӈ���h���ƭ�刪t0�G9�դ(Z�&� br�\ۨP�J�ÚdɆ�aQ����d��	"bB�@\�ĉxNH?t��p��q�����.^]��
�.e�DF1D�C��ĝA[���I=�|��T��Tcmd�<�Ȃ��8I>H ��H�5l;wڲeKS2��9>�>%�c�N���xO[k��z�h��֬Y㩤}2A��[���ݞ"@�Cؤ���B���ǟ�} o��4vh<��U��0kĖ����u�9��4�6a����k.�-"[��SSS���c�/AZ������W�E6�ţ�~�����7V�̹�Jl�h0��(s_M�����<��*����{����0��J��2)�!�]@���.���!f���}�h߭����� �F+$D�%Z\*�W�Z��JaJi�z�*M�	9
p)d�A+Di��Spm* ���l���YbH)����BJV�l��3�3q4;�V����1;y�$d����y���}�݇g���9�{|hH��3
6*򁛼���F���rȄ�3�D$S.W�
��OaVԁ�=O�"�/6��xG"ϟ�+z)��4�w6��S��q#LB(ɪ�j��R�)�P�VxXi��`�<��JTX��KB\�%b����2R+��Je2�^f�x9�Jy�������4�A�^R�uG��P�x0�ь���C���`Ӿ�/ם�m�V��{���t���Ш�~�ee�:Tt��b�Br<��C���Lzff*�E#�����ɜ�bYL�����;n�Rөn,Y�0��f�F�81�U� �䳻�&`V�
���
5ye���*�&eDS,Ab�Xh�BT�~���Q�����t(]��q�/��dC�[�������r�3��)2��N�Z�A��z�'/�)�%jN�)��Ҕ�L�C�;4g� R�L�"4��R�^�6ٰ��ѩU�q���؄ÎD�A-h��eP�<!�3_���/܎�Dle)###�I(�z�h#��	V���4��#27�QH�<��B���s���;�E���F�\q� ��H�ȰX�y���&�%��5LR�Cj+�^����5y2�ʅ���~<���U��:(N�J�X�B5�S��3sx�dD�^��!^�/"\Q�s�f�������u��@�J���;�H�R�$E���#��2�<�3�.�[A���G��aDOEܥ8>�mTJ��]�J��4�&��ǹ�+��Ǐ�h�n������ɭ!��I�2�>�+X�p�����q|	v�c�`.�.�ɴ�8��'z8���Ygi��2L���dK��GI�����w�<752��_��e�`��޽{I'�ō7vt�$׿��o����χ�:D6'H)�f�$�=����w�;9t�[nimK�!�c�p�
YJ��I��8��1�*r��ל��m�Rfs4�OSC��"��|a�Z�t�.���y*AL�
u���	sDX,��X��'����
*�2�{�' B#���x.u6�X�aժU���$����3.�������NGW'��|�f0&�p�'O��S/]F�bp��,��	�W`�ES4F��QΜ9��d�Q�2���M��݃����j�~���¸7�=K4�h���)k �mJ�۰��N���~-����	\�����8o�Bæ�e��b<I1��ޑ�M�R8�,Y���{'��s���4��о#�������~����4�і=�v�F|��p��`y�1gQ�~&#@�&�Z"zf��t��X�WX�"� tE��O�jעևH:̱���d"�e��G����jqeBY����u������x}S��?zI�;h��Ԯ�	w��;𯳓F(:����c�����[�n���6����L&�����
Lj�t�nG"4"&���VӴ���ڻ��=�V�,��0עBwvr���ڻښ[�q37������C��9��h��}����`2���œ�{T�՟�̧���;�g��oh��#�Gx �˖�Y�����"4�<M�u-��̓O��¡��E۶ި#��m�4G��ѕ���=C*�Ы֨���4Z�dފ�h��MI�p��^�Ixԙ�<�O�VCrp�a	�S�;J��MA����ĮZKߕH�3���tI��Ҫ�[�����p��]���\�W(������پ��	��[�k�y�MU)��υ}��ሐ��OPjM��<�⵷�˪D)�b��9�L��Dn�7=�7L*����r<�\��!����E�q����R�5!z/�;RS�9� �e�%;�/P���%8��n"���4���NNbB��CΦ&�P�~�TJ�,H8՚�%g�G(&�z{�@���{Q�m���S?��߸��ŋNM��Wnx�(������n��vFennv��t��Z��L���UkA��N��x,��0�/4�2�F��>57��GN���}>ͯ�O�Jr'�>��\nN�����q���Y�9.�Hf��7-x�i���0���H2w���{�NM�t�9۷.X�`zz�a�\�)�,�kW]u�5�\�/}i`����pd�]�������Τ~��C+��̔�UVx���׾v"�G�!�&r���5Q�3ܾ��o��׿�H����ܼU�MM�ksG��Z�#�N:��QK5�FN��,�m޲���QW���$Q�+(�ӧOGB�ts�`�"���Ä.^�B�N��+�9-���&�!|z�V����cu?�VE���^Dٓ(�Ň]�i��]ԏO��2S$b�e������K��m#���ZA�
�G`mhE�=\���J3�X�F������;=���*Pg%B���(xb�����(I���H�,8�%�, 
R_�JQ�� E������(��6��˺��Q������v}�y�	�$kױ&�K�K�5��T������5I�_RT��1�K���*?1�<��5�e��E[�l���To�)�1x�>�����<���#!�$FYB��P0�]��҄VQx�����/����������𤄺
E�F"8���/T�Z����8'��e)ލy6�_*�Μ:ӵ��sWo'�Tn�>_���/�	�3y�Z����X��A�?�<��h�
�KI����c�v��?y�<I�6F�̌/Gx���f�~���t�MU��gϞ��q�� ]���e����Z�ﳷ��M����ۭU�k����3sǗ��ggZ;:����q���.蹯|�˸���}�X�k>�b�&J��V�sV�Z52vl��1�#`D#٦�K��tEPB����w�l��ݒ�=��#�ٕ���.Kp,�����Jh�l��xz����Z
Q�唎9���=�ܓc'�\��4��$%n����*�^�)��D�o[T��x��x�m��-��M��ZQ�`��֖�h���Y��i���xAȥ��?HcU<���/��B��LOC��%¬B�q���a'��sl��VO�*֌O�OQ��UI��a14��rD�f��נH�	QRdh��;��s%�*����͏LSc�I)k������Gu�X�@�l���J����mD��x��i��`f�ahj��d�k�ܒb�����uJA8��IHr4t�`��`�|Yac�j�V}:Z��l)�''O���k֬��=��������ӡ�g���+G�X�[����˯N����|	.�'>���?����S���EKs���z�Rƃ6��@��A�����˗���\z�e�S��P����⊫�=��!��_x(�ϦM�p*ZZ24��OE��[ZN�i�+����ۏ���Z9�I$�"U#D6��v�!�^��+�m���/�ʅÇ���B���
N�.]����/���k�+��@<U%����QN�#�������η�651��Ҝ����DF?1=Nԉ��T`'C$���e�z,���	��/-�V)�x�IFNCY<��,T��A��R��1=��u&A�b}�$��� �i{��_��V����7��_�R���
�.��,�2�I�4�
v�ïe�ܲ$;��1��R��h��x�c0�Y���׈��������E �[E��0��DzwS�(�g�ă)�������X�@.M�B�#������BǗJ��\�9?��TJ�NIZ$�%�QO�V��Ls�~��"�JE���5�����<�*=r�h,
�@���ge��a���K�dy���D��4p.�HR�e3��.���@�H�lM''˨�b�����PYZ�R}!J!+pYq�[[; f�gFi��NL�Aʕy���o�(��iJP߃&K8]�6�������(�4���D65;sW����S��n�z��6�d,�Dx>��O���*\%p�f.�!���a�n��c��?v�7��꫸1L���$�4���M�x�	è�^�n���,���[�w�]����/�����/�ǈ��z�����X<y�M�j��B�O1�m\����MQ,�uW���d����B���[�&�M��������G׬Y}�eW<��#�%�81 q������sI0�Z������BI�J�V��gN�7�p�}r�rMj0,;^�����)(�z�lG[��,�ϭ
i��ޕ"Ľ=F�y�:�i�0W��i�Z��('F[��&"���k4j�#`�� ��c-b�:�y��`����v�
.�
�J�A{�x�S(�`:�!��Ō2쪹�?7��$��J�4���}��v�Z���0]٦����*E�!f=�n�ć>v�e��_���D�.�a�^w�TJ�q���+��(�.��j��kk#V=4�����k�B0��axy���ilCZ�l�"{��WM�7�c��\�"C�F��qr�ְlA�ES�&?k�jН��+�,�[*F8�\!�
�*jƱ����2[�5rP4����E\���4:&@)��Q������2��Ɋz���v�K$���1�w�i<�ݨ;N]V�d5(�OE�����b7[���t�%�v��#�r|ZCM����[�b���#�/�̧����}��A�x��^ҿ���)x����w86>9=3��N�߿'��M��'��k�m��7�p��ԙ���V����������¤��ڎ;<�����A��(���+��~��w�!�'?��w�}w盯�ќ4�a�l�
b0�Sw�y��`W�;����侷�s��Cp�9�C�*8�]1���ܾ};�>�QjǷO�%�c$�c1>3�+$��и�%`3jrɗ�#�Vɏ7JDs�Ra3B�V�(�.�8���0:KX	�L411ٷ��%;�� y��d���XE�^*a�f'�hSY߯�t{��PO��vh��K�;����e�/PK����sLe	ǨT�B��q��b���b������#k)8ա�!՗�f�:��,X�ןɟaTd3�������!�B�5�A"1�|�$�5"Y��(�X��/�D�>%<,Ҁ"Bp�F���X�qiz�4;�ݜf8[�̨?IΤ���MN��sBV�M�xB ��C�)�
�S])�73>/ ����B�`tA���,ã�IS�XezE
p>�Bɠ��Q�y&Cy��4c�&�RGW��+�qp_qo�x��t���5M%8v�á$k���5g���"����~��OQ�l�q^��f����ļ��p⊅�c!B���#�k�s�N�2l ������Ͽ随��}�^�0A8ذ��O·�Eȃ#@�,���g�h8�Ϛ�vզH�5��gBV�������+/�2�H|����ۻ��֩:�JԱ:�����7\�훶o{�{��	�����y�2-��������i?�w3q�k��޿kߙ���k7a����u�R�`$�D�Xl67�l�1a��kT̪'�=>�b{�����bͬ�s5*�)���,��Ru��(x�	8n�V�u��X U�P$S-�k}C@���ɵ`�{z!rݒ5MUJC�F���#�����eF�߻�~8�L���UfY?��I9��~�?6�3����%)j��H�	�v3Ĳ\���hj�s�����T�0<���zu�QTM������5XUz:���Q-"�
�֠��f��=�PRfk�0�޴�3���w2�d:���YNˢ�8ʵ�#A���sqSnݠj��Q�W��Y%���#���j��ko�V���p�`�Բ�N����v���1��z)�3Ê kB�^놧e��JP�����K�	on"0z��P�q&��*�Q�JB�`ͫEx�6�	
 Wj�e��pL���F=�(�u���Zɨ��?;[��#7nٲEM$��_��Ө��Z�"*p^5E��N�\1���� 3W]���g����O�<��R�*$Q�.,S�i�mCծ[���	b���E�z��?a��?���2�+a��Zvb"ߞ�vl���Kϝҭ핺���C�[��j# �G�x4^�ϾQ&B�pB�8�	5::�bŊ��{����~��������]G�}k��˖-{�v��Vs[��uU�����x�	�����+:9(gll�7�rWO� eHb[[[��v�Mƒ���!6Q��0~ N���&��%�J�(��T!����s���ԣ(�T���Bn~nF<�����T�iY�_��װ�v����S��Z2�D� 	��i��{����zb?�яBIR�G	8LA=�����������s�{o��&��V��e��м��N9LS<��e|���_�79N�<!^x��ӧ֯_/������b=5cѦ�����*�"T�'��0�iW���2Y��ea�s�ph�y�}F`#���?$�*F�.]:R����D�l�������[�v�X�w�:N�޽{O쟇5�� �ѱc�8p�탕7��m)>J���а-a"�*�M��;���j��_����a J��?��?\~�yX���3U�`�Ƨ�C�-[������{�֛�ŉmq`��8��5�Q/�c�XG٨Q��˜���SQJL�M�-*����Z�j׫/�����7qOPdJjbC�����ے!,�w��"
�#���z���!�xO8�I��,�ƍ�.]�;����/<��]��g���o����1*�r��D��f��$���j��ÿǳ��}z�$�p����ή�L
"��f]�I$R�l~.K3ʛ��
���̗j�>�#��=�f����H�^���w�/+0��L&���Qc��Yw����8X�笉�'�na�8&�n��ƚHW�y��L�-�i$�F�ٔ-�hx�*��Trī�jB,T+:#`��%����Q� Dմs�<M�4O�N��=]�ǧ���ڕ��A�Y������%ч�;DE�&�I����c�O;����/��T��o����,��]�:�+�X*,N��?%c�2��������ߦ:�L(���c�;w��������MO�y��ֲk�|U���D{ �0j9��-�;98�/ώ��-\�fb~���k��d�z ;T�hskw��k}�W[ZZ�Z�lq��M]v�9#��a��,�~�
y!�zVk[f��:=<4O��3�𩫮ޔnM.�Z�w�'%ݪ�}M��J�%�N�K���F��h ��z��>��^�V���jZ�*s��o��d����$x�Si�ř_<��n\Җ	�M��Dp�ь��k����&�5�����Z�)z��ʮW��"�E�惌9a�}�uT�RS��g9�d�ԝ#�A�ԋZЫW�T*���N��T*��|x��{9�T�R#�8�ڶ9cH<���?��'��̝߀�}�ϳLL��\v�����zp6�&& �cc�����]>!L%38�-;���65e�6�B<�6��沥��f� PQ[�̘D�p�|�`x�%H�7���X��w�@ ��-����������ԧ>OD���5����s�E�(��h$�h�l��漳1:�����(ԘϘ�ȮJDk�m�Z��ț�9��
J�{&{uΪF�Ae���ӲX��Xߖ�9&���,cyi��ye���6>	���,Z��V*����������1~{j'��6<2���7�(x��ɓPuGN���+����z4��܊�n��w�y� ��L�6B�5/a3\)�ʳY�№�O9������a��e���V�OeJa��O���Ѧ,i4AF�(p��ԩS8=�FR��s##Ͽ������*�����7�Q���̉���5k.\�������~�f]}����ba�;���nݺui�E�kp/��BG�,bƦ#!�Ha#�}ĳ��-�2���RY���]�r卉��!�L'-G��4wZp���=�NԲY�SKx|Φ�c"�[Zf�
As-���F�(�ě�Q�h��+%���5��9W��=�/�ʀ(���!���?���
 M��'�|���׍���9{t�y�A%�c��E,��c���B�2j����a?;��Ks�s�
�/tn�(��X��_adkk��?Q��W�]��_�j>���������e��ax�ذ��L��N�r���Ǟ=!OB�'�Z�<s�7�h�l��_��P���/�}���KK�,y��g���_���F��LF֬Z\�O4Eԡb����f�*�D��m�y�@hg��5����R�k�E����FUr-��؛x���i�]��'_(�#��ꑰ�G@B��4���*���gR�bM�˪�����ó���>}xa���O~�;��$���%�׺�Q��T-<��Yb�����Z��;w���}wz۹��h����8<�IO-�ڂC|�`Œ���D˒k��8�hUQ�W������wl3��>|8���?����{�n>l5v�4$Zz�fJ���ѨO�����DǪ�x$ݲ�k�=��*z}�`g�~/y��r�('���w�Tgdyɒ�7%O�|;�%����I���[Ӳ|��2\��_���Y�E���\�]���X~���pD�o��hh�"��5��O�9>����e�W<�;Z�Ѳ��dV_��kn����/�|�T1[�p����G����~����Z��lh�_E��F����N�u��k ��d�ʫ��]
4$�g�F^��p(ب�Y�
v)ն�T_W��
�%c��
I��P�m�4�C/ĒK�@gU�o���F����L�� �J��-
�)MTB�ٞOT��󹂠�:��j�qzfp���������ٗ��Roo�@����G��^�Y��	���Vb��n�y[o�ozЙ���JP��-�J�k ��V�(��~@\��?���>����`��c-Z䚤�z{/^�iEm�=t��&	�V�B��[izp� ��5/���O�l?�a�G?��_��Ц�(լ�-{��#�֪Uk֬z뭷�q����?���Mص�5z�A�\?)�r��	E�����y�e���~�k_{��gz�!W�5���Ztd:��Y%�X��q��;C�w�°Q/��g�ʕ��0Dp��9���~����w���р�~���=tz����Ͽ�!.�R�1pl��#G`O�q�g�y����*���M{�UqD���uH/���^��̨]�Vh�=S���y`t��'�8c;�G�����
�h�B���y����r������M�C<>�ξ}���*� y
���_|���/�$�����D���SOam/��R(&ǥ��W\�iӦF��~�C'��4��?���Wނ�u��^�l������yǯ�ر���?6v�����]z�������x֥�c��|�M6�#
%>_!HS���h8��2��\�O��X�'�����c.K�N�%�:���c}DNf
��g�Ga���(����T��R8;(���IYT�P>)�p����6���6�ă�bU/M"�1``>[��5���&�S����4%۰'��p��W@@fgw��t;Ivv6LGU���I<QшsF��k �"�����`K{۹睃u߿wowGׇ>���L�u��t���l��I~��/J�7o,�ʜ�qX��c���-�����S��MXr�Uc���a�Q���{m�A�c�tX�����i�lQ�c�Il$E�Yt�cCn<�~�G�\>��;�8N�5q�
ցf��)"�)=���{���ǧ����l۶�[��.��`7gRD�����������?z��M���l��/���[��7�h2��������O�Q����/��ʵۄP�����hKk�Өb�%U�͖�����r�}������-�=�jB�Ν�׬����Q1j�W�����g��_S�8'����A.M^7Z�!8=1�����o�y흶6x�����'�����##�m��r����՟���/=�fkk�}�%��_�m׮]�s�sp��e-ͭ��X���)�|�c;=0�ё��e8H7�ݽ{�+�<~bvӦ���6G-^l�{�ǿ�{U{W��7_����kX�8�3b�6
+^W�מ�cI+ʲe��p��c���h�D(خ�Q���������-M��Cn_��k+��=yfX֏�y���@0ܚ�5��;���I�-ٓ��X����=P���o���/���k��hk���/bI����榦��*7�H�S��rnzd&�W)=
�����!\x��m�Hh���#�Rb�8b<�U�z�a�^
������o���*Ň��tmERΏ ���#�SI����A��UN���&d_���) ĺҽ}=�P����}Źlehd��Ф�	�Pl���@�:��L��|#B;,�sO?}��ю��qEQ��?�!�ْ%�8i7q���@m��W_	����C�I��wp��k׬�����#�q���nD�M�0�mTg�_<*�Dw��mx�X�����K�N�~
��/kt�����J3|�Ƒz�{����b��4I7�� =����ݳ����Dx�wt$e�1 �*����q�_s��'�|��j�P���矻�ٷ�W_}����/���ŋ`͒�à�w���盆�_���򹅟��s����aq Z�_~9q��h�Ÿ�i<�?��SS�8E	�V.CI�"=��7����O]}��د�	�&�o\��P%�M����981;��,j�b^y��A]I�6�Q�K�ň��|ŪTE���ɦ$�`L�ܔNc�C>ײ����l��-�8�Gd�x4\��c�߯��(�G�Lu��c�?������{���x�TS�aA0p�x�}���3��޵W�����7���D�D�r�=��}����߼1$�V���>��O~��{�X��+�2��Pܭ����h����9#�	1�a��hD-�H�K�8�D����.��5>IC]i�\�
+Ɠ��05����o�vގ�o�ytb����۷o�h�y8{'����[�nn~nL,��c#�ՊY7<�v�FS4|���{���_��u�|4�nٲ9���l,v��~��[���X�,;@�8�PQ�?��?~����o���K5,�C�_������7�1t>�'?b'�=�y�M�.���Q�0V������z=�-	��f�&�E�Ѩ��3  >��~1�i_�r��;��_T�>2:Y3힅}o����M� ��iDR\�RY�fS��P����dl��ǆ��������o��,�bq�bQT⩵m��F��j:���*�X���E��}�L"F,ƆI�BrP�)������?�:�w��П�
.Z��ƕ6��_�*4KG��P�.��5k��o��-\�q3u<k�#DX*#�����b����\�Pq�ݲ{��N�M�t4w��F}ާ�ِ�$�7�;�rjh��u���zc�+���n������4@N$[�F0l~��iu���K�eǕUI�M
Z �۷d�{G2����EF=|��d*�8��޳��P������P�Ͷ��R��c�u+��kϷ��D�ԩ(���ٳ�w���}���t�T�5�M����������Y%�^ꖠڒ�[7l�t������8����788p ��y����'>h��=�$fr��hP/���F�m;w�lN�|�n���̹�b"�uճm���n'�NI��;���7�~��p�G�>?�}9477��Y8<�����pÕ*a�O�<��$��ݑ����p4b5� #��㶶����Ȼ_]��sK�mA̕I)�`#�k�a�#����)���;o�>�=>t��Z�����z���3^��;$�o���-��r�UW-Y�����NPGYs&��/ 4�������D�0]���iƓ>|���n�����B�~�������������?|����)/�4X;������?+7������i6�5C�Ƒ��6)mX�U�ޙ�r�'����_���>��:�$��D\d�a3ƴ�\6�Zᗳ1�ʑ#���j8�_��W�kV���Y�v�N-��O�#�\r�����Yai���9�8�7Mi�����DF��{O`��D��xŕ�U"���Ћ����	�Y�c�=�ܺu���bKK�>�[��Z[F��	ш"�	y8(#�m�`n�̧�"��4	��[��֎s.��{�}��"A�k�3���8N����;�/^xp߾'N@q�ؔ�kW���9Dة�ɹu떘��n� 5�JH��NK&M����._�c���YRdD;X�W_}VoƚE��JG���}�I~�+�<#�d�ad^~�e�n��
���-�cx��S��0��`ς^���J��Nо�Z�h)VL�ig�8G#��"Me�N�J�M�����E����zR�eϢiSø�i�|T�a܂�z�i4N�}0�p��f��-Ɏ�����~�'��[����a�qw�,ߞO�HQ��d<n;��O>�ܓOc�r�yʧ,�+H}&S16�1GtF6�m`�|lt0���4)�<22���<�\�#��a���q����`8!Z�W*UN�:�K�'�>~��cQ5_�ĉ�����&`���2�f�5	�}'��w#Ѧ'�zRd\���(��H$���~,�K��{����@�Ju>�S��5��U+�����tʗ�����{���_��G�I��Fc�H4��ގ�C��|�[_��y睴2'i�=��{qkG�����Ew�˄l���}�/[��[5l�����W]�x���+V�^M��'Oa=O�sfhh��ձ����MU�zKO{0��-�/5��Jyxج���cA�A؞��d�~���R�����\s|BJQD�z�"������������#W�^=����^�̭�n����?$�-[Ⱥ�\�����B�dM���7��?�g�������\���cYS3�>��j��p����/��N$��xcjjjrn�)������V
F���*+����B%��7BJG'��F�X�E��j�Q{Z�ͷ�����8uz��»ẏj�Lɚި������>[�io�>B� Mb0�tSPg
�A��۲�/�'��.7�'?3����g�:p`K�H�A�Ό���CWЀZѽz�:;_P}b<�D�ؑ��V���#��s��}1����'���yghr�3X$��Ru�QK�XS8|�er�,�fٌ�q�ف��+�v����G��ⴭvG�&��]ǂV*e(?(�j�
G���穐�/��톢ad���Ƚ�<�� 4�ta����KY�G�zKs�a�ñ�8N$�u���C=��@0T�a���V9g��p
�}��Te����aA��~�/ϴ4�LMC�^��"�z�ac�&a:��1[Z�"#>8r���+xy�2�V����F�MV�}F��������]|��0_%�D��Y��m���rՄڂ������w�G>�KDYP�Am���ݩ�>�V�R;&M��Ⱙ�8���po,[�$���v����vZ�` ��BR�M\
��?�����۱z�����T��S����A�{m���?/���u�]tZt*�il~�����c��K����ߗ���i��9VԬ���ڼ}�Q�GFF ��W!�|JYGGҪ�5��x���虳�N���q)���w��a�&�s�q�:&�,��B�!]��d�l�ʹ�q�)�vƶf1�&ء��G�ylx,�L��r�!�q��;YԷO]���pB�A��v����t�1@�Fɏ�\���>����u��rت��C���YR�?�&91fr�Cn6j�b�1�R�G�A������c
�����юk�>ITj�*��D��0�.y���+����RK��̼���3�L4�ע�,��OM�T5h[��(*�
�U73"�sYqc�H#�ML�f2�Z���Ȳa֭����~Msi��_3����\A��:eg�v���Z��ӟ����?lڼ��O߸{�[�G���^s=D��
�A�&��%����7S���I�*�XS�VOśq�f��2��啦s98��욙����C��b�ߌC�4���4`��H3���ɾ�T"m��3>/�ı�fn����6�;�oaw�N�J5O�ά[�n��߾��GG�Gǆ�uA�V*%xe�Qv��_{G�;{�����w�9���ts*���KO��Zֺ>�Wg�����DL���ο��:}�0�C
b{:VT�����)b��Ս�Y.%�J�>:|�>4x4� �:F�j  ��IDAT#����S�?����l�ѩ�֬Ye�汣Ǟ{�u�����? �x�jw>xhê�VI�I�ha�I����sY�<Y���W�"2�i�>��a�U�P�r\�lӵݢQPd��%RG%��i4$��X$��!G���Ir�,�3�X���j�1/A9���c��Oƛx�8й4���mVY����yĺ4�HLS���'h�`$��e5lfK8����"!'�v��W>�J|�T��?'�\c��i��E�T�.��P��mrA%j�FM4u�!Q�k!�mm�i�&��*�����&;t��S��٠X.�/�����'��IU�dL��P�f��W.]����:�X�3V�p�����A�I%���՜8��Y���������o�?E�8Ma������]]]�]ǡ���K`L�!b�Y'��Z�B���<����]z饰��~\���Ӗ������FS��O|�=��K���麨/yz�-FJ�*��Al{GJd3w᰹������o`�>z�ex�C���iƫ(�Z��!����8��I�4'���m�V�<���e?��L�HR`��c�3͸�L2�aÆ7�yJ�Ǉ��ƭ"���L�do���'��I�1���٘$��'��^F�y��A,�z	��!�Ӹ�t[�e+T>��s�r*4N?{��珏P�oc/���)��6Z'B�e0��MԂ!f$�<�P�h���m3�t����8)\�
�M�R4j[+V����ܿc-�4�ŵ��Q/K�(���i:�\Y��I��$vb^��eAV��'�ٹ�l���	D�ˍT�_��O�e3��y	N89E.�>��Z�R�)�����
����yt|
�@��aٔ5��9�^�mۖx,��Q- (Ky�|������%�T*6�r���4Pmq5�|�����Y�ڶ�3��5�!�~���>�����#�k�`K
Q
�g$�ؾy{a����S_����Y�_Ũb!����k�X���t��L�@T����Ӭ����q��R}|,;>:�t��d<eV�$А����xSK����o~jN�|�lX�(��4�b��ɉ�QS܆&'Ϝ�_�lJ�f:�� ��Q�ss���֎T8El��	�p�Ё���ݯ�*�\zQwg�k�
N_�O��hF�i˰O�ɴ%�-5L�F]u��������"�T%���B��f�&�?b�Z����5/�Eî��[ګ�E�����(��j�<YZ�r��;uj�gr*���MM�`�2)�a5��ۖp��Qg$�䓅t"
�)�V��y�ꦣ���Q�$dyy��,��iT��|��o~�>�>x ]����¥��08~&�
E��~��p	#��Ǐ���������*��t�V]�tn��0^`�Mגʥ�?�'vpFn/�D��ѹ�1c`�=�bE7 ڞ��LH��e�'�:A��5��Hnk��h�E��geV�h��I9�ș�L�AF>$ot�ީ������!�t���(w'��e3�m6���d���Ɖ������`�%V���BI�[3��o�1��b���"����A<�ܸq#��b����g36+���f<��><��v�@��C�ǎ:�8q����N�V��9�;i���ķ@��W�Odc9x�z䧧a�"M��<�&�H�נr󄌁1���X��O������"���Suq�P7P��jT����!6r���#`��X��[�f;>c����yFA
��[��%�%D����Z��N$�%ϡy��?���D� ɦ ��)�l$ķන�]�V9����]���M7݄`��bYԣ ���4|B]��NQ�As3K;_��O��2���%�W1���2����hj��E�~�Dٰn-�YǬ*�+W�<a�%FyǞ[��˖@��m�"	,>⤤.���coIDA$�l�b	�������EO�Sk���~"���E6��nV�?V��I̶�f��;�bE�,7�h}*q�	ĳ�"��>�nҰ&�n������!*o2�ǆq���
qZ��T��X`CI�Ӭ�=��1|���?q|٠2F���9�2�mX�/�Uk׭��jm�Ƶ�p�ٛyꩧbz����������%x��_B�l���F�6�a�qMF%YO�v�ф��Z�{���7���;l��q5��*�~���\D���%����qV��k���M���ok'�BDŲ�kin[���ٰ�X�`�)_�F�1����d+&f#�@󦭧�F�z�]�V�e-b��8�4�fT��;N��_r�Ѡ�H"�.�nmxlT���s�C�]�qI��gq2�nފ�loY�Օ��R�LeR��a$���DS̨�����6���ݻ������7Mɂ��i�g�ZR]�i�w	�$FIQu�@p*7���Z�ٴPEܺ�\�Q
��^x�k6n����Vj��'�H�����5�����d2ޒi���4u��4���W|����������lO44��"���N�Nڐ&:rv�|zh4�-�����П>5@��%=��F��t�kbe�� ���wށS�hYhp�#Ӕv����Q%���2����;k�ۧ�݌����<�l��,h�ʧ��ʩ�䤨��ϋ�d�,�#�1�&_��Ţ���	�d�y�<���R/����)�$A����Nv��{s��;�z�� cM�d��ҹ1al�Y�EBCs���]pj��$bU���+<�����6^u�n��n�$�}���¹�d%;9�z ����9�1:�d�i&0�Ƶ�컗^}Ib�E��"�o�=Ku�}��� T�����p�\9v����i���V��,���P0����Y���矇�{��}=��M�������{��U��ç�s����df�$��	]Y]�UQDQԏ\��]�Etٕuumk�EiR%!�IH�L2��;��S���<眹a��'Μ9������|�N�U#6�1�uEYf��{�lK��KQ��b����r���o[9k���_��p�xZ�v}�/�P[׹�g�}ۂ�kli�%ٳ�20�z�%�\�[`+�|��3G�ʭA�ѧ�zjzf]�b��w�=6:����#��v���Od֦I�^ҋW��S������r:;U�~����L��?�������G���K����{n4޼�EX����s�^l��.E	R�.��Ukz7n�(�u��	D^G�ug}%sPH�F��tx".N'� ��v�����:�DX���c�{=��V�>�CW\��&���(�M�P�87��,�+��>	b`E܀�����S�ؼ`��w4�L@��s��а�#A���-���	K�R)[���J?G5�rUF�1`NbIjv�h�ٔ��wu��+��:�6�� ���LN�r�9�|�4��Q�1p�ß �Л;5ݞ��tP�&��������>x|��էƣ��L�����F	6rTU��EM�����dFW��rs��3�2 Ԧ�[v}��"C�Jf�¯!Z?� �bs��k����������`��y�ʒ���n�v�M��Mgf�f����_&��5���i_һ������	�z������8w���^)+�d���.�+VA�S��2�X<Z��[�����+��|�?�c)FY�#�X���o'VO����縪?�~���?��\{ƅ���m�O�>r�ʸ�J:���f���l��~r�� ���֝`9t|���r�
��M�#e����O_�fg@��֮�Oe*`�7��b�"}݉Li���Sٶs������#�|���������(\�aÓ]=��(�W������~�Xӄ�-���7�=�H1�����\�Z �e�3~�I� ���QΡbj�XJ���6B�c��cWg��E�'��<�W`���!3[,��::D���V'�&���+W��#6�6{P��?I�}���vW%��@��o�Em�G5h3��gE�dXB�b}4�Sᙔ�Yq'm@���8]8��K-�3"F<�Fme�r���Y�����%���
F"TO]�0��j�fɐJ��]���bP�c����{�"O��T8Ӝ�Jb4��a�M����R�#s<|��f�ٹ) �buN��A����_�oL�я~439�����߻����~�0Yb+V�X{�y�]C�cT��8d*N
Y�
*q@4I��T��ԥ+C�J� �:��"�%0Rۂ ��z��Jy�uL��b�9��K_KWWH�������K�((�b�7�Ә��d{z�I�M�R��A��FnXR���U�"��Q����q}���o�X�lM>�(fh�m,�Z��D1p��K�F�� �LnWXP�T�f��Ց+xǎT7`8�]��:j<��O.(n�_,SӪ�_~yff6YO�JHoii)��/�í�hFWc�s�M�ⓝ���<� ���$�fNO��&Z����j$�v�&M\�oh�t��i�,5���d�%8H�~t*;�S;�xl�AV�[���Ȩ�!Yv�����)e�J��T]3d=}אEM�૊g�
t�P���%��֒�8Vxd2p�N�S뜰XX����V�l��6�4gEq"죆~r�r�<v2�����(� f�ms��8��&g&�#ѽ�:�����{z�ڻ:��ob�.W�<U�4�3�N�%1Ф�jut���,&�p$��hB;5߆��W�l$F��]�l�G!+r��T,F6�6�N�%n�ȕ�.�D�|&����AI���}�7o^�r�7��k���}����EKV��M���Pk:��y�E\ڲ�(�("��B>�0ϸ���L�@�xϣ3E3�[[�"&uζ�PMM<6y�&,G�ćDh�N��n̎�H�'Rqn�umŮ:4�5�Z�3QWW_��d�?�j�'��],�hČiܕ���+�I5�Y�i�[nN��|5oh��̄CD(OQ.ȲU+(I=KN#=�M �5=�-�2��±z	y����jluh�Q6���d&)V�L�[�R�T�\8J��T���J�:Q�/���Y8J�����@S�9�h�����^\�!.vM��M��nb�O�:��\>�iF1�3ʺ�&�Q�T��'ca�����HW�� �=����G�F�N�T���Zȓw���Τy*V$�#F��ml��3!f��kT�FF�j,�ƚ����dt�e6�CF���������ۛ[&'�#�� O�(��IE��'����LĔa���j�p�����޴�I�M��i�BN��b�cH�l61�|�r���f�[�o{��7����'OaR��IM�KŪ����'�;:B�\f���ފ㙙
;���Uq(�/(����d���דּ΢�:%I���[ܤ��\�wIF�޽�W|W��f$LC���Ώ���3A2��e���ߏ�wr�\���	�͸p���-k�Lt
�X?��$�#)�%�6WLI���'đ
���@���[�����a1��
�x���
q�a�Q�s=wp�n7�YD�����aU�io�Fb9":M��d8�t����RdA9  m�'xL�H�����$'� �1�|.�	nQ�ٽ�6 ��ңH���<ҙ42�\��%9�%���o�n��\��� |D���'ȏ�T�t�\��Fym`��T���y�6�����Cm��Ƹ�X���5E��+ �jm�塸� �Ek�׹�9���ѣ�l���o�$�uʒ�h2$N�Ax8�Ns�yMa��2�ް�O9���R��	�Dr� ץ��(s�H?X���8	�5'���$�_r�m۶m|n����3s��;x�`2/�+��i(�r�248|��'�����0�c�Q��:��ᡑ��fq�0�%LZ,�H@��ࡲe�LN�p�l&Wu�$��Ԙ alh{s�r��W9����;��h82p�Ϟ=�-��S�ܥ4�Ii��#��E"�r���U���E�t߾V|۠j[�r)��T��FA�l�*����I������\2n5Ǡ�w�->� �%�^Ѹ��m�e�Z�w�W�W�d�%�琸���%�,>-a��al�.��(�����d.vo��<����x���s��<�����R�^��2�=�aVm�;��Lp�2��PNY#y�A����{h�@�,�e����f}�^�Lφ������0H�)O�-��ֻ���+�8[^}����.�RHk�7�D!lN�/ҽ���X��&'3]�}4L"��>�t�+ C�U)W��V���1'�,�8�]�z���,�kA;ͷ�¸���~��� ^�l3lP��c���
-)�`f������]S� ݬ���<���'>�|�rn�3ۺu���~�}��U�<��Ï��jk��s�4"ۀ�n����m�v|��O�ڵ+����:��{�����|���mx�5��[VV�
��R��׾�5�j��?v�ʕ����C�
s��@(89&"S-����#|X�i8v����/��#���3*W͒�Ub!R���"�D"�v��U�;�&$�c���E�'�	���\��0�K5��F&˞%H(�b�%�xi��	F�ќ�9��@%кU��3L��źT��珐��i�HV�.�&ĺ����ɢ�M���2�W��<D	�
m��I��]���r��<^��a�)H��[�� D�1�ys�4	ɱ���(x��9)/KT1�i���%�g��-��}饗�}�Y�Kn��q���GB�6�tLNO84��l�|�H�P	�!�[����Kv�ų7#l��r��U�B��Zu�iw}���^ziNQ��?��o|�3��̇?t3��׿���~��lv����Y�E�k�N;��kN�ڋEK `�]��T������OnٲL�Ԕ��J�R�VxL��qa�+_���SOݷoߦ-���NC�$SсcG����u�]�m]w�q�⥋n��\&[N�#QS�\MJ�\?r�  ��׭[�w��ڵ�O~}���������ɏۖS������Zkk�T&
�ڤ1��(�*�Z;�4IZe�V���-S��L!�����ASW�W7��u˖��>�#<f`+��0c(.��(V"^���Ѓ�u-�F������j�,��*{Du�[��Ad]5�ƅ�ɭ/EMq���CB���y�8�q`(�G�\�l3�hg�����ꒄr��g���R��OԱ�,33#ߢ4	W��{���`tUA����o�P�YsɫG#���(�-MT%g�4�-�w��a"�B,cv�u*�'�T(и�Pk�(��oR&�<��w���c��K��y���4�\qr�9W�b�ؿ��?��@�5l?ޟND�G3�y��I�:��#K�*���m���-��S�q^�M3�F XB
E�����}���@зT��7����o�����'?�g��_��g4G�XH�✔��\ur���+V���~��g�q��ŋ�[{c�N��-�k�s�o�� �G{[7�0XF��xqBi����S3�͛7���kÁ��_yha������{߿lٲk�������o���461��E1 ���g�[�uL���+��iO_�����c�}��W^y�O>�����(&hP���"�i4W���⋒�������u4��K�}�Bo�"9TF���Bu<�6������S��,�;�	Iz�^H��x!fZ��[+A.ţ��8uA�� CGqE�Rf��,�@*Y��\\p+�����/1Ӛ��m�Ok9��L�1Ye��c�$�f���*GY�J����,$-`iA�^�Ds�
��R����K<��RC%P,&4�k�&�p2M*M5V��Knp q5-!ʍ���ZT��#1�pI�����5�fe�3y �+o�r\�GRI�$����!�$ ��I���v�aA��5K�U��&���x�G�3����w�wS�@�����/}�+PK{橏}�c��ݯH��5��Ngu�H\�~�����~���d��ܵgc�=��=��v��-Չ ҄��EJߴA'�����>M��ƨ[���W�k��ՓS�P��XX�o��&(��SV����������K)����v�\�~z����w|��-[_��[�����s��:;�@44"d�"��].��3#�p�R�?~{oD����f�e>뼵�V=?&,�b����d�`xĀ�Hs���R�(R���*����|�=L�H-��j� �!g[�o�j���Z*M�S��r�V
f�劬���0�l��|�y�4����k�cĴ�H���9eQ��b�_����r>'����!٩�19��b����~E�'�c�&��+���!	��&yDz�a���>�����PS��L_ojJ&c��[hT��Bْ��?s�M_��|��y!����E���z�r��U����
.Q-ނeG��;��5�5Z;:��G�ɔbs.�ư�Ƣ�p(LXײ���&�i����H0��PS��ӱ�I�=��݀�c��i��`���X<̋�)��?�^\�����u`��O>yph�С#�&��S�V�����7mٲy+컏~�ݑDtْ��O:�嗎W�)3�mB���LOC�-\���]o�4�c.�#���.]L]>�)Kp.G`��[o}�ǨvC�\�<55%{�������|��7>��/v�mŊ�X졇���������l�����/�u�}o���)�����&��Z{;�\�tuSEU��ӡu 5�T���K.�M�կ~�&�'h"B2M���RYB�B��	�|�&zHi�7W9K�NhG)���$"���HKR���iD��*F�dc��$ B}�-IMx�LN����q��j�<A�3B@ނ`e>��rr�p��G���U�HqY���aϡ.����cLs�S���L�oI�
��l#�Al�sM�N�we��+K�ǟ�Z�p/?���VGFFn��m����ͯ@H�{iT���(��u�?4o�
ϫM�zʙ��B����Ν;���Bs6�m"�`�Ep	
J�2{��꒳|�A-A#J˜�|�=��\��H8�p#��v��Q
Mgp�%K��S�2�G�#G��ÇC�www_����K@�Pร!���.�#�cC�#ؽ�X2�ry�X6!�Gc]��,�.�{�gէ��l��Z,M2�Nر�>������7�ػha4�����O|���$2�ҏح(�� l__���OY���Fy!c���/]�d��U�Ja��A����f�,�sC]���/���/��P����
1_t�HP��@��u����S���\	Q޻V��XbNE��	�KPK>���f�!�6X,������3��l�q��)[U��A�\��u4
���J�H>!�F#^l�	y�κ��&ʖxV��Q��<��T��6��:8�"ǥ磙YQ����fk�y�P�^����)T�� @ǰ�
@�ք9�׵y X��0<���̮^�-�1��E���|��H,�y���)�CN�hgFF�]'t�W]rɥ�p|�֭N�@o͢^G�2�Y���ƪ�O�w�ҥ���abs5bj��C��v^S��G��T+����+��lfN�:�����?�Q��ə�G�˭���}��7����7��tC���Λ\�-�������k掝;{���=}ݫ�'Y��\�����]Yߴx(��:7�A,H ������v�9Cπ��o�����꫸�9k���s"����)K���}���{�}O<�DcK6����s�=w�U���|����t���k��!�^��x�t}*���������v�J]o�:�$q?��N�AQq�#��bK�,�hk���@�¦ݸq#�������]�@�h��aKd��U/j'�0A�d:5�U��)��z�F�U�+��K����;���~�"��U�0��:�xwĕ�lV����<@|t#O��JE�)��4P�D��Z3���r�8?�L�,Ѩ��Mn���_s@+Q�[K�Q~U�_����F$��@5re�HS��<�_AH����EE�9.��1*��h}���K�1/8��[/
��`��p_K;�Hf�T�Z.GSa� ��sm|��(C?gsg磏>�۔��P��/��W�ٶm�W^)�
�ۢ�4���zN,C%�����f�zD�L� 0*Т](@UN��A����ٓ���:T>U")B3���B��Xg��wtte2s�b�#�^x�f �x!l+33;t|��zb�hrm,�z≧���߇c�E������ܲ���BM���N�������ax�N.W0�4�`�ʜ@�߇��uM�u�&��YQӓ3
c�6�D��������?�яnڴill���#A Ʌ>,Yd��٪�)(���m+ J�+$��ԙU��'���7C��V5����x�ȠR��5�7)�"�Fr��r*V�#W,��$R�I2��b��U�L�
d*er<��4P��s�,a?�D;(�>�iKqUՑ":���.P��/�-Hu�|KP�p/��)�ɜ�5Y�#�}��� X�b9r0�D�FX7���OLN~���7�q�}�I�J�$���g������~` �0�mD#��;v]y��{�\�X��^l��c���qh�	�+o����_��ҝ���S��ͤ�h�]��ɤʖ:�� @�|BW�46R.aQ��zk��闿��/~�k �H�f0�-�r�l�&(?���M���ѱ��ɩ�斆B%�鵗w��s>�<Mե�Z�+��43o�2(\F�<�������޷_�Zг�زe� ��S�tR�&M����aФ�Jew�}������nuu��]�uXef���C���hnw��FO��U���"
�=�1��fMe���R���A��3�{�$<9N������-�t���\K�')n+n���;��Q2�'�A��Ӕ?��R,��.k� 4G/�Zr&�Ggn��X`쑍�y=(��0�x�+��[��Ľ!ZN~�I쵫��خ_T �gQ�8a@
�]w��\P��L�-��gm�i^��吅&�DQ����[�d"$��=]Me��Ǹ�XƮԧ��x�|���>�005ʭ4���i:N���E��|��VQ�P��K�?�H��j���+b{�0��t�\eF�J^�)�?�tӍ���6��iL%w�ƿPwب�����!v��-�ܲ����<�̵�]mU�BfR�8��+�RC8��B�(b;�fཡ�!<�)�onj��+90���!�������E���ޡ��p$r뭷�-����?���040p�EW}�s�,3�h���!nn��-[����W�X�8�ؔ�2���ѷ��T�-V
���x�#g�:�X2�L�f�>��+VAΥ�)���瞆�a��YR�p/�������	lKg�#�D�CͰ�GȆ^�&�5H��}�t�Fzy4�
c	�	W�J�#VR)�H4VG.�S��Һ�.�8�蜰����b��\q���FB9��ث�	���6uCW\��pi� ]d�����D�/'�:�$����(\��{�\����*�sAamM��B<`/�1�к��(�s����J`��T����V�F���j�!�"6%�ð/�_��C��puhnG�45��9�(�S�]С�v�\��	nܰa��ŋO?��R����ut4T�v"�bGT��ѣј�����5bl@�J٘���X3����cy�r�R�œ��o~��o��ƅ�C�u���)*[(�����e�����/>?]�Z�f�t������Zw)	�p�63YT%��4hB��c�^&����?��;�M* �M�^�=�40�������I�����u ܄3!�	�PpA_��2�C!� b��gi�֧o�����4ա�`C A}0��b�9���]�Q�N�@-&8659>h��@��vV�����{�<
WR)ǟU+�QPU���{S��S?A`3Y:�X���_-z��Z��U+"��D��Xĉoyj�5���X�(�>R��Ur������yב��>� �R�e%��&�g��՚�9����=���%�F��'x�q��U?y@�7�l�@aC����S.Kgjj`|�u'qi	9J�\DT:�P��޸F�F2}�SJ�]�(q�����xӨ(Y�<�v�v�a�1���n��u���qS��!���%\���fU֭[w��k@-�J�,MQW����w��ݱh{�sKE�Pe1x.�3W�{�������g^|��_[/_���.��D�w����-'��*��!������ڵ��Y�@�?��?c�^z�E�Ժ����,� ���/�B�{���h<�ĥR	�Shpp�uх����ݪ��뮅��8p�ʳ.��I���Fc�B	��r� s:-���J�fN��G�tD�b�"6��rV�
u�u���s֞~��.��ד�]��ұH43��Z��l�R%�ZuQ!#�*��L�`�F�Z\reښ�Z���,���m�'��Q��t��#�c:{D%t�,A^LC�&����lW����TZr@O���%�/�)����^�����eʊ� b��h]"�������!v������ZkS�2��r���,+�jM?(\��.K��<5�(b���'8�e) B�
��)��z٭�7�+�Rf�@��9���re�hS.�U�T����-��c�Peֲ����#;�Z��B32�WĠ����|��׽�R2$b$b��!HV;y.A�dU	��rs���j.��.J���pV{{��3OŞ��<��	�<6���m��g(�w���%������?��O>�,[�lpp���r�)X�3^8�����6��C)Da��Ѓx}�����ʕ+-곥���=��a�$[,˶��v� �����hW(YJ��$Iǉ)��mR �䪎G)f��L���t�N�#�E�$H8��ǋ/򜵭�lV�]���~a�@���F~3��{��!��D%Z���U�[��ɩ�9�OHmQ������9�����RQ�A^x��	�{��e%��y,�"��(Ƽ��O0BJ�7U��,X�?�����-��TM����Bxk�ý�b��uq2�v��h��"�V�G*���|Y��|+�e�%��ؘ�y��D�Z�;�g�����P�mp>�X�O��U-r� 9� �l�)�Ln�*f:���/���bb"��#�C�F��Q(B)�W]u%40�\6]���C�3�p�N8�w]��I�%�J�J� ѷ�~�駟��U�`)�(�C-��B������7�?�ɿ�p�\pA4�e&{.�K�U�[_���o}k��[V._���
�*���&~�P���7���+_|����fH�K���1��ͨ��ёi�5K�)��*69��9�ډE�'����7�V��O^��G����=܅�\5�b��:�b��:����b�ӏ���0ê�3��B��� A1õL��|(]�X~� ~"#�yR���H���-��!�*��0�%tOr^� 3����b!����+#�Y�&�\%�9XM#2#PX���V��"q�h��d�V-�'B
�I�ɪ)���r�8�X�\�6�{$tH�)~��#���N[�I��U��9#-9}�Wa6J}a���L�Η��q�lP_�fO+�_���,�7�0��ũ���?�jE�rU����+�b��c㥹�%�
Ź#��?��>��bh��ƆOL�<���J��Phlf���Hܰ��X�j��-[1���ܔ�V�}�����������?|{�n��F�HѪ@O\���,]�XaӬ��T'`�].����3?�'���  Z�����LՂ&{v��[{*�ub��eZ5�P�v�'hS`��x��{�h�����T]U��sP�/=�<�Y�|1M�9v���)�cccؾ��:k��/�q�?��ϻ�;��^Z���~�Z��ZS�^ޔ	��&�����uv�����8�	��䓖�����[��xk�ѵ#G�P (ɤ�	��`�)ر f��Em�B���(�ap���-nި�1��T>AP^�I�m�3a9qr���+��"�^��l��I��m^J;�u�L�ќ����;G����P��`=��j��t��~e`pMQt�)��{�R:2�'5�U��vׁJ�f(%��!ŵK��\*�N�����GT���C�hf)V1�9���w�����}v��������(y�#���a0!Xn�ҥ�?�SX��Lߒ:LF���5>>i.�����'�A�H�0���8������я~mD�[�����0����C۷o7�!)g�=)��4��[�m۶`5�w������]�z�]�ׯ}$457�M!�eBZC�J{%Ibğ�c�2%F�a�%Z�-x�|)o�*����L6G3�$P1==�j�I�C�/�肖�&\mxb;���5����3\������yS�]�K	���\�d	Hmٲ�`��>����HGw5��M
`��S���B�b����Ԫ�Lv��9��BfW����"a�/�j�1%�'�h�"5(�<�T�`}-��ťBF�qm���B��f��D���|����'R��AЗ�^�  t�\�P�ӫ�՘�՚�I _��+:/,'�Q�5���c!q\�&e-T���g`z�g5/�H>�a��Ij�|%�Q�o��&X^��S|s@�[c���֧>�������x2A�w�j�a�65��L��ܷo-��(��ChW-Q�î05q����e�"�x�9T�}�D(Է����ף�>�Db����H�5��M�p#(��R�H��?ө��,���uo��s�MS;�s�)J4?��Xn��o�ٳ�V�qsU1�%6-M;�V��>��ދq�Z6��]���EZ�לh���cs�9awy���[
^%��Z�Cm��-^֢�_2Y��X�y a #�4�������}`#��z8 �Z�7�\���%��8�87��ܚ
�"GlB�n�� (�*؉��W�?��Rk�ɧbU�"
X�����(J�����'��{��7���J�!�#��㧧��7TӉV�R
++�_3�{5���6݀���TW�}H��?���شkZz�U�J��Nb��(�dr*5�r<T|[T�1�/����V��(�������%�%P9�JU+e�Lc}�a[�h�HU�r��?&��Hf�J�\jP�:<4$����b�����YBQ�/�l��ݷ�p��'��L�D�x���;��V�^�NiWZ�ɛ���4�^xI�@��},��Bq�ש(\ �����<��t��W��lǣQ�����㢣K�ʩ����723���FJ��jS��n�i������!��ϷuPc��T[����-��dc��b���R���82�
��|�J����HD~0�GN��$fR~��2�f�
'" ��T�ڮ��Gr߈��jK7��������h�30���'���:/�����+T?KF�S[?�O��:G�B��+���@�����-���u$yJ���,�#Bܢ������9T
�K��KƕVS����i�j�Ȥ\S�K{a�$���kW!� wŇ�A�K��y����yi1�	ʼV�[^C0Q��5��d3�L�x4���׻��w��{v���dkk{OOdv6}5>9�P�H�ʯ¡��"�b$���4峳�A�-
��0�q98xd��E#�9�_F�T��/Z�Gk+WLݨ��Z�|���115�����D$L=�b��(�����=��:�C�o�����
����j�A��{k�$�yT��8��(�R�gQ&5%���ƯbҐ�7��U*	�$)��>	S���cO��+VlX�?���[��\�&?�\VJ,�k$ˍ(��T�tQ�ů|a����T;UQ$)�JF#M���^B	U��㟚x��wY�]pk�r�׀D|�(Y/^h��H\�V#Y`�%D	W���%(�T�Ex��>Gl*#��������y�쒥)O'��W���#�W��t���Z����N�� ,�+�+$İ������VO��,3�I��I�K�ٙ���?�t�M���pc_O7M�l����N����&nGD�T�Y)�K	*�L��{���ϒ��Fi�B9�EIcY[4J%����쵦��M�6��yі�d&H�P��_P��3s\���n%�ϕJ��U˜d�� 
J.���p�zȶ���]�����54Ҭ�<e͑�I$����)0!��|.�+ԥb�ExwX�5ف*U��I�ݬr$�fPd,�(��5:�R_�f͙g����&:.STЪ��8�(���oE�`g��޺u��*�J�q��x����fg2ԋ��I�
�+v�m��wO�C0[���xA��p�E�)����tL�����$4i�>`l9@*�����("��_#U&hS�9&�\�:P��"U��� ![��<����&�x�у�'6\�hK8/��Z�l�"ɕdw�i0���A��	d��\��CN�
�4vC��=�3G�OZ���.�BA�U��W�:���{�IO��mnHS�����מ�j�����K@�S���B�4ƿ����jF(�c�޽G�i'O%�l�B!U_�z�:7gPg3yy��x�j�Jɮ�V._���su�+6L�J�Z.iIMN��9�|�˛�T�3`7$�T�2����R�"�[�=xrJU�
ZQ\f$A(<D���d���
=Ğ:��@�_���@ْ�'��d����zQW�V�f���q��<����Ӝ���c�~��_��?.Z����g���W�6$������ķR2λ�,,B|v�}%�����5�	D�ԟZ��d`�Gb���C!
:�ʖ��HA��Cb��W�TF�2���0���`�Y�֔}��)��A?��rq�[����A���3����q��%y�ݿu���rN��zՃ��W:8��duځ�	���N�@4�I۫@F��B>G���s_Dr���	��(��F�8�Xe9�� @,-�J�nA��-�<1T*��b�SD�]��-�L��svxɌH���Ef粁Z��,T�2�1%���$�=+<����)�;p��,b��;K�}Ja����0�`��.]�-G��x&�qʎd!��7V>;ǂ/��p���0KJ��٢:iJU����M�sHC��MMԂ)����U+���" �ŉ�1��#n�њ�ݻw�V+�k�Ii�Yg��~���I�Ymm@�x�ɑ<�F�Ú�4����`�,�ԣ� ���qK���Qj�b����T G�$�Vtis̛����ڳ��(
.�j��}S��T���H��W�`����k��X86���Q*�r"8�
D�������m�{�/$��#AzM�㪰�����܃�UU���A6��zXw������Ё�2�.]/���G�"������ƙ�C���PBtC�Z!�`S�'��Q3�F���SuҐ1����z	�WAѥ"�vU���
�9�](Ec��?
 �5��
�j���&��Z��s$uO�X�n(���q���qDR��McS���JJJ��CD��=o�؊�%c��b�
�jC�rS�Tx:�)��p��fi�juU+V��D���D���硢�)��%��J74���p����Sg\y啯n�!�/|�ΝbB���wR� ���7��mt?q�Rzi��PM91J�6���P�0`p��mg>N��F&S��O/��{�GUko���Yܚ4No�;?^(O��k�#|��"�QP�-$���	>�g�&�r?i�v��i5E'�Sp�|�w��~F����+܋��	(�A�0mH�T]��j�*H^в��EP���dGGGss�F����q��Ύ��G��'q��@Ҽ4���ڼ����� ��-HgJ�i��e⇮�'�b2��4��L���؁1/�X�-�o���aY`D�.�������D,�~8��	X��+)\^��j�"������?V�DC*�w�TxT�K��io�,���YD��/��k)A���'W���gMǆUX��ӓ�����w���p͝o��;��b��C��@���<��#x4l+t��8 �H�K~kײ/ e:�'D�����SK��8➐��D��>�t�'P`z�GjM�m`Y�~zo�Ew��,d�bb��H�&~�ʿ�xGk��p4U��B�\����;N'%�gu.H'���ٺ��W���(��&��+��))g>,!/H��$ �%�R?���I��e2RZ�#C�NªX�E���h̻��/8���Ѯ����F�rSSK}S#H�T����9��	tnm	�a�]��+2XHq�N݁3��i��p��\�zb�\/9I������m,G�j��㉢�+��!I!'��=<f�!�������9�j�T*G�j�R�IǓ�7QUDjR3�rB!j�o(Ӹ��U��RjKZ�"��9u�d��=s�9[$�9~�;���<۲e��+�>�̋y�Qöm۰�X��� T���n
˶�����sk�yB�~��g �K�>1�&�3���A��k �Ф���<�p��0	}Qsko�3�"v�S�vDC*'�`��UN�̟P�������"/]��&�(X��<^o�|����鬪�Q�s����e����qؗ#*A�R�� �i�2�͗a�_�`ql�(�D��R�]M�LԲ�ͷ@�-Mu�ǽT��8~���c��.�X�ɤ^p�/|	��
^9ԉ(�V���}\+l�)�7,��1�@'���,�i N���F�jBW�t��'�J��fs ��9 sG�Pc5�ؿ� ��S8���Jc�]�\��p\"KH���Z�h�K/�41=C�>U��>Y�O�jܚ�	��]��fX��Ñ�}��+��bB��VҪ Q��s�nDM�gfzzz���w���y�w�`[˻q�U+��߿bl|G�P�R�υ`:�kW-�X��EĎ�	H�k����<4{�>F�!^Y�*9�B�D�De@H��(�������q�_(��v���k�P+,Ti���E��=~P4,%��5���HC GܚFX�]�)�\p��r�R���#oUP��&$�X"�,�yԢQX%�!��4��Pz2/���������%馦�Z�������V[#�\�Dqi��k�G'0��(�C�>����,�`�p$<��8�j0���Q�;@�d"-A�|�
&+6��lR���:��4̻��@�;r����:�6���K���5k�<������Q|a.�]�~��CG���-�
�������!�0<r�з�����������Zq2���������[?q�5�\��k��B ��Vl2U.��6�{������ ����Mu8xph߾}u����0�Lv�F�[�n�5�5�R4OoxZW��n�Lܪ]R}�#`?��i����� "�Ц{bX�������)�LhH��
y����	��;x����ϣ_)�1Z��j)\� m�R}@�_?J!}�,�����ޞ�;����8X�ȁ�?��m������9|"����O��-`cQ)�+,�J�Y)-�{{iT���4N�b�4�钋>��8���@?��2wY��ƣ�K��u@ϳs�8�dmd��}O%�kd�\t���9��X6G��5.*���h<��kl{[����(�o�禄i$�i"R�\q��#��u�}�b���~�?��d2>22�������-ڴy����w�����l��4O����I���r1-^�d�ƍ�_��o����Dp�W���\�w4�qa�I�ȨE�_?6�������kcas˦W�o���/�c�+V`��⾫oh�ϸ6���������\q=��+/=w�}��?�v*�2áB1o�F���t-$	G�p}_B�tc@dB|��eB�D'�r��o���X��j���i5U]Ή�y�+�p>��g���0�"�%v >�]��i�w�Fp?gu>UEV�� �:A�^�3��AN�m�����Z�aǸ�c��\�������`Ϊ�}TAV��?��b�Fs���2=���f)b�XO=����n���r�Yg�˥����C�����N�8]�
p�<CfhtD7��ʖ��rMgɋ[ߊ�W��iS�R�H:�+��Efi5���D���-��v��]����\��Z@;rlp���[^}���^�Z
8b6[��k֜J��B'���A�|�3������~��c����$��]�s�9�o��?��W_���C-�ĸ�B�+�i�&�.pz_oߓO>�:�m������߅�UW��$ƥ�t]�Zi3L����<���^������'�|�o�[�Jd>�-mؔ|���3���;���d�dL]}΄a��S���Wy��[	����N��ꢖjߡ坆V`��Dɺ��GL�0c͠za���2����ݥ&���X�KIu汱�k�Ԯ�%�~E�����]�֭�r!J�^�~Ϩ��[�4���4������'^�.@~���,%M���S!�T�Oj^�"�У�>��o9�&I*۲eK:e�oذ�V�M�68No\58&�#�E�	���A�E�n]�DR�/�����t�b��<z��rr����t%Y\�Ġ���!����w�E�x�����B�U�<�u�駟q��_v�������������u�I'Q�l���%U�����k�w���o~�<XW[;88���[��Q9�E�]u�m������
�}���7�ʅ�먉HX���u�H�x��u�u��g� L�%�UOŒq� 먐/�v�ėl}b,�J2�����_���N�չ��\�ů|vl�����O�� ?��RU�o���O@U���$C�4H#Z�ho/�OV�Jes.���9p�^�+���`q��t�H^�t�ג��ڒ�^�.��聳��!P�8���ĐS��G�ܤF��q�p#(��y�Bxl����e�א�4n &|\�~�}�h G����6w	� V�"��8~཰��[�I����.�x=�z��	%�!�|T�͐��B���i���T�PI�[Uu����� �%>Js7U��`;U�hאNEg���i�E�;�:�55j~cCv��OL�n�|�l[#���[�'3Sm�z�Y�������ב��lmU$i3����2�6ν«Qw+N~6g�C���C��J}G���D[���''�
�k����(�+I3T�NOM���H,�'�-����e�?u�m`�]�w�?���Q*�6/^����o|��{���{���O?��p�P�����%���"A��@�K�.}��g_y�@�z K�ŦAD��.�蒉T��知��t�$D�^��V�����_�����;�����Ʈ�<��G���s��$�;k�f(�r��V-_q���Dr�Q#��۷bU��O�����}����X�j�پ��]�X�D�:�T��o�o��D��~U%&y}��8�!.� "*V�҂��S<-*ՀA��@;����E�1 �Q�[8�y�2��sbxMV(DY�3���C�t�?��è������wީ��Q��rBz�5+\�BIԛ�[���j ��b.�\��괇�&�*�T z�W��g���a#�5<��f��cy���O�z��+�x�':���Z�����o�43
ƞ�/����ݺ�h0�E�izS��rC����%�U��y�@��cIx�%�֮���ƒ��\�!>l��"���'����m�m��tu�`��Ũƿ)i�uw���=|��}����lX�r$澀�X�}ջ.���m۶-\���k��5�F����z˭Z���w�zsjr<m_����o����oq��;�HW#�
S�����?��?~���=e�I��\q��;�0+N�0���(�=g�-����X�|�۷n��f23�����${ͻ��رchh���w�i��hi�t�	����TK178Lc�`�ON6G��j�[�K�v�9�{*��t���N�	c<7@��ϴBX|&��W"=�E����DH&�@�o��Lr�Kkֈ�mWR����,�Ƴ2/D���k���6��Ae�;��̀?�@��4�9��)�p\?�K":$P�<5��[C,dW�5���&v�;X��0DW��*b�
�C�S��m�۩�k�[Pn���MM744�|���B���|l��w�:12fj��&X��ÙY��LSJI"^�8L��Z�O��u�1h�9W)�$�mN���J[j5j�������h[[��W_�gϛ@���X}S����Ͻ��t���ߵk����YN;��j��"{����h\�LQc�x�u��׿������cc��i�;Q�b���XW������ ���)������Y�`A��3�̩���q^u�\��[`��~�}vj�+_��G`b\�=�_X�)d& ����!8�OS�Q~x��|�;˗-}���>���?ץ����
��ɑ���.�=}@��9
-�9?ۑ
P��7���J�K,���O����|��ҹ�G���4�4YBhZ�7��T��nL���{
J<�� � .���o�����Z��_��滧�+ीs�V�g�y6��g�a�uj0�� �)��""qBt������v)O��$����9�~B5��S<��{^/3��3Z%2�Ȉ�eJY�WRHֻ��N�|�_��W�:6>J;p���:��t��x�cK��y�~���DW7�XT��&��o~wij�A�iܗ��
?s�t뭷�~�Y��	W�����﯃ր9������������r7 ��	��~�c�z���������뭝[6�v�i�Z!Y4
��7J�����ЁDU���2�cbtoo���B��7��b�����g׻v�[)��R�%��cQ�=��**�Ҳ�+�����W�:v���U���C��ݻ��m�J�/w���4���T����!>%�Ք)���Z�)�4��<�LN>�T�zȮ�b�+!��������w��}�g�u�-Y�d��C��X}�5������Ur��8�\@$zM�?��a�]"
�	k	�F�HdL��R2��NQCT鋿H�S�g�
�"g����1;+O`<͏ SP��|/<�?�O;����0y�R�a�Ձ��S6oL�p��G��=��)�V��	�"Mȝ(����0Pי�$�N���.�}ⵢ��t�JUI}b��N�ȧ�&� �*��P4a|�&�R�홂eFR��'�!j�;��uB�MQ!
���Es���(�\J�0�|���S�����)sǙs��{�}��K/��׾>=v|ѲE��:�����^ݥW\���ͷV�Ze�z")~ho���!���K�hj視vgbr�q�p�13���O�.<��ӵL &��8�7�+�a����Ẻ: �څ=��R����-5�� ������P������7��r<�z��o��Fh�|.�m�}��{�Q�{�R3�L&G��L3(�jllZ�h��%u�oS�m��#��ٖ���h�z�Id�������X���]Yu������H�ide�RrBT�R�N�R̶��YB�{R b��{]���)L3���wk<��ΩIuEۋ�)�$�����7f��RP~]sf�Q��8��G;��>`�Z&����%���5��@~`�I]����$�q�/h�֏���q,��Ԁa�Ւ%/�x �~>�n�ԑ[Px�D�{zz@���8�0;9'b�rD��>mV)O��г�,.X�܌��Ž����ֆ�����q;%\u�2�yՕI5w�u���>�����t�u�}��_����{e�d�`��L��8D�7�͈8�	}}}˖-,<�K%r�qƏ�E0�C`��Vh�5t�f�������q��;_=>��~��?�]{&p}�0������4�;<:|�Yg�~�mXb$������E��c��>������
��y��]��Ꚋ���Tjhd�Ҋ
����L��MNOK�P�/n<��3���� ���Y�|y�Bm!q����4��i;ӫ�s��I�k�����>��Ƽ�<�X�?���dv��yU4!�پ��C2��� bR5.�`\��k�%&^KP�N��ەrG�� B�����0�J������B�@��kJ9�8Tj<@ Z����)���3"&Ƴ��\����.sb�ns�ꅵ覼N�~�+�Q��"�hY�T��>�墷Z��[����Xn�XQ*E*��I��Ü�f@E�cXR[K������T�cO<�r���N_�{n�K�|n6��`��EXF�z
�U?wG�~���c�ܜV/��2H����w�ř���?���o������w�L����-^�8z|0��>���R�uɐ�T��|����ƺ(L��s��!jiD#nx>���n�,��M��s���/~��s��ݳ����͑	S#	�QqT�ܼy3����G��N˽�#7��z��! ���o���[�_q�%�z���߿�3[(�p&'��;9fgg�Z+V��ԧSt#C��%��>%e��Ҧ'�ݻwr��z*�D�=~�x2a�i��"JE��8S��Gj��<�
B.�����@	�#��څ��!zBxG����2x�(,���.W����Y]���爩�	�ﮯ(��ml���:�Qkݚj=�/&�h�(��e"�T�I�}���X�
W��� �jq�U]�t�`�*':��LIי*�'��q�h�1�Kğ��,�>U�4�SInv�_43�;����@ɢ--��� *j@��FI7JAa���K@T�H���ѣG�zϻ��_���hf,#�U�������冟�0�T����꫅�Q�|�ȑ���/~�v��E)v����(L�T(F����䫛7'�ug�u�������ͯ�s�9�>p�yg�%�N��3@� pX%��# ��sY)H�).�K_�҆@�߻�[�x6. ċ/=�ӟ���gsjOZ-t��CG�M�T���%��F����q�F���ÖUI%1B�6�4^t�Ыǎ����M0|̌A������)�nݺu;6��E�j�RC.�5���Z��r�	lH��q�F �ٕr;׏�C*PK���xIj";uv'����/�cy�D�܍Wê��eV���hk��|V�	t�s�VK�̤|8Ҩyi7�ϓ��AAi�K��A~j4�R���r";�a���J�F�Kf^���RW��Q�P$
��?��������y����!����e�����d�p���FdW�����=5z���\A�`�k~��ɑ�T*�ixff�/~Lx�9���n��uǎװ�u�x"\�,�\�jonn��db�v��4���D���\](g���n�����N�	�q�#�<��}(
&��р�]�R/=��G��F,�07���[v���Vjq���4�_/;M�h:�ɺu�|����d���r�)�΢9]�\.���z������z�ɠ'�K�!IA��7���;�'�馛T�� �tuu-Y��7�hh�s��<�a���*uL��/�b�?Bd2{�{���O<�4ͩܷo_c�}ٲe�b���B	���/Ǝ;��MI�c�Jy!!B KY0v ����@���</�����:~��Ց�x��rP�䭍rI��9">�U�SG@����R�Wgr�R�6��x'7�����?��Z3o0PSb�Q���+�����3%���ѼA~�*G8�}�(�MF�A,L�<.&�2>��E���$�,L�Y�:a��F��/]R��]ݱhReH�����,y�MͫG�J \�z`���ڽ{��W_��/�m�wH��\.�S(T�	� ��{Hc�*3��#{����v�W�"M&�#�E�+n�]�0yQ��4�rҼ���Sߦ|~�J3��όǁl��T��趓���lk?r�@�삞'�|���g�������ȑ�W\yUgWGSs���s����sll�\������������\>]ӳoA�Kh	�s�yن����@����T���޾.��B)O���15>8!z��IT:�3L&P�7��~�[}���}����8/�С~Xۛ6m:s�Jr$�S�l�[����1�{�ڃ>�rR��'�b���Մ�Uͥ6��	&�;?i^�(5 i��C����5���:��q��␠T�#o6O��|^��QR� ��}�������	��j|?n�Xr}��M�aN��D~�}(\'����9�Ȯ����:���p�x�CRhKV:GS�!rG�M4�����+�.�F�D�B�0�G�U��T�LǣԂ<�/�
SS\dg�Mh�����O}��Gzz�+���ڙg�m�괜jcsScS�l&1Q��xg4/�T�j����fS�E97�Yhk�"��5776�e���������I��|�O��'�{��ϒN�928QW�N�E���Fw��65v�'�1�U������~���~����7�|3VI���ncA�|��MLL�=g-�P" &�\\a���?����rfj:��M�R���u���>�WKA�jY|B��t2-&_�B��[o�|���'|eѢEx�p,.���㧬X��)A��0�^���]����:;� ��)� ��Ui�#�����3!�&&&pZ?_QLA7�X�~:yK�msu?C���8���{4�̑��OŅ${S�5�Oȴ,ǝO�����L��:��Nݙ�޴��E��^%�ݴ q  �bJ�b�I�˟%!BIBB�8��c��.�EV�Vm%m������=��;Ϸ�?�ٙ;����w�{���駿4RΌE{��}1��4���ä�(LHϴ�jB�d38L��9��a����SDz�N�D�#q���>A���i���0A#��$·�#W� {�j�z�O��Px�8*n��bŊb_:��N����=W�Z������b�L8[�n�C�Eʪ�e�Ru)�1SV�@����#%&��S�Q,�v:\�"R��pVj�TR#�P�+@f���826>77a޲e���2ȪҜ��^��b����q|�ՓO>�{��n�	u��t�������ʕ�k���P��m6�9�g-�h���|�;�q}�-[�7n�99{��a����J��������prV���	z��g~���S+������������D��(ގ �p۰ux��������ݨcwrYJIܷ7�y��{�?���?�X�
�/$�K�ǐI��^�~UGU�F����$sT,ԭ�ݫt�Ie\�Cx,j��EM�v:n��\�Mw�3/���t��_殖�R_�1p�f�0�?�����9y��%'�t�� �F����s��[r@:O��$:�b��^2��.�O��݋���r6a��'Ӕ��Q�i��5*�o'X4#UA�'H7���'�ŷ��� 8��
� ���)�t�����'e�}�Feit��2��C�����ݱc���(�sHCG<xb�j�C�_}��
�b������/���#��"�U����mwt�5��bB3�nv�^@]�b�+kg��P����c�]xbinfq�t���o}�p(n��Vxd��\m��8vtia~�]x���o�n�:ŴU���-�����&B4,�����3�l��e�����ڵ�>N���2�i8���H����_�l���@E��~��D��P3ccR�'6�|f�b�DU8Wz�\�� �%.u�=���)~�"ɥ���_���$b2�����iT�2��T��m������7�,���Ӥ�֯:e���靽�t�D[$:d�c�R�"�V\�W$����G;��wf�(HK?!�Q�F��m���gm[��N�\��������rN�8,��d�Y�3��K����2�%
�|B���#��q�%l�F¤�#�:���XJ0,�{�\4�q��&*�G�#��Rd�vy2W&�+���lc�ݞ�C[���~ �"C�O�� !m��7�5�_X������G�T�O[�u��xˍ8��s�V+�^�qb��h��1͠dLˡ�p�G��dv�J4K��L-��X�._�\��!~6l�\��Ү7`��9�n��εkW��!`�cC�t)�2ȱ��A��.�Q�٬7�D�_�8�?{}Z���9'~俰};l&ք�GOH�:izt�y�V����H��y��4��_���5�'��ǏCu���ivo��}0k؛_��ׯ���w��s��U�O���OZڗ���S&�H�(dw�M���ͭ�E���(I#��9�{��%��0 ���fS1�Ԍ�@K|9����=�,9cn��ù�\������t+:��9MZ��)\A��*Dή��x���݊
_�14i4�r�'Go�xO�6���A��;�d�T��éUxr���ʐ���>�����t>Jo�QᲪ�B>d�6O���
�%x��G����\��@�&����p/l��ͲwCMgl��f���k�sLS��9}e�$q���*UM
��#���F^7����|����X�0A��\X����^~N���7ih�����x��V��Si7`�&pO�=3�l����i��Q
��mu��\ffv�Ӧ�����C�f&'mY03�N�9�`�f����f#���zj��ِ臚>��	��W-I�K}�ã�O�+���'��;�ĉ]�b9�S�,��P��/&g����f�3�gH�&�������R�Fq��)���L���/�g��q�]tQi��霬��/A#XF+R��_"N�J��KQQh�o���=��R#�fD��X���d4<(�,Re�G�R��+�}I�.f)"��s�Ak#�I�R)Bs{VW��|�� �0��A?�5| -�F8��=�򜜘I�҄�ǵ�ũ&ߌ;%�Q!�ɞ9��^	G�Y�%A-!t�O��J�E�C	����#��.��k��_��/��k׮���7�:vl���P�xR3G�U����o9p����w�E_�
q���hj&K�"������@U�����fu}�� �j���r�F�2�*d��/-,���<��"uW �h�hK���� ]�2���$,2�^���j=�RbR�"l��p��Yby.�Z�Ӏ�a3s4w�7S1(��qCJ1h�`�[�âDz�6��Wk-��)���'���Sk�B����KuȔm)K���������i���T*m�e��w[���i���`v����B����5Ÿ�?�긙��Ě]a224qأ	ƒ��\&�Q���nE
��y�`�<f����X@��ә�&��.�8�/'E�����H3��h
ȨxR٣]���ɤ�8�?��0@@�9P��C���W���H�#Cڱ�J�4��w��e��#J�d(���3���a�cm�abr[���'e���"�=�25οG�v���$|M�/��jJL�:nʶ�n̛J��O��h�N�w����F�g����b>�I�E��6T���)�v��~���4GX�g�:��:��0�C���%��N�@T��o����/E��/�%.`��v�I��jE�l>��z��c뚫��L`xЃJ�5u-�h���d�L�m�J��N�l�s�(�C9���㜩
�M���1��ڗ&]�yVZ;>{2S���#�x���=?X�z*)��8c�7$j:�u�-x�m���F
�]8͒��{�<R�M$�p$�����lJJ#�Lco^b	A<IVf�K���p;��`Q�����*�v��S�i�O�l��-��Eׯϕ9����A�~�	�JKc��c�A?	)���R��Z̤?'1�N�T���Ҁ~-���-�,�a��i�NV�C	W�p�5i.����5��e1�Q@�A�����17M��ٮt�KD��T��Ȥ�7���66�F�ʊU�te�q�;��?*���vez��%"2�P&Ր��)���u�\0d奫� gl�y"0�r�O-����h�������JS�V���P�q�'�:i���%`e���S��0:��D�N��=Ay��F�Y��o@2ߗ�ù�$��ȑ#۶m{��'#?��d�{�'Z2���mK��K���}j��)H���bBU&�������y���$�F�O��=�P^��2ɨ*4���i��G;�J�#�r)� �b�©4R܀T�aФ%��\���f2KLn@2x*���C�JS
�P|G=A�S0�.0
>���[i�Q�}�Jsq��
h)�Mw�'H̈�B��+���ByQ�_R��*ر,|� ����o'
N3�8n�`K��͢&&5Y	cAe��?2	�a6�u�q���_*�#���>�cB��1��!>C�fy'�
y1p(��Yv)�Q�.G�ְT&�l�/�7l{�.u�em:E�}YRB�&�*��Vv�� 7�?�h��p5��V�VÝb#�_|��'w��9:>6>>���]x�ʵ+sC�����Y0-g�1CY/�%(<J]ƽ`��x�=� �d��INH�:�V/�+��ƦҨ����b�Os�'L��˩������J��E�Y�|r��Uh�Sb�x��g����Nە� �i�Ф�r]�サx20��na�KeR�C��*B��O$6���pGIO��;4�C(���-��z��-q���\�l�spp!l�|LF�_N�n��|6���5C���U��&���Q׹C�&}�G��gr�S�o��/��#��R���jc��n0?

k����s�+���D��0j�zqr�C}޽(�Ɛ	��驩���r�v8��H����H����L�
 ���t�h: 	�W�Az��HRa��\����wdm$�Gw&�M��Q��V�Ғohhzʈ�7�@z~��#n�R�EI�pbb"c�����<��S�TvժU�F��^�2�իWw��'�SCܞ��	�gt�n�1�������+G.C{��v�wb�j�|�O�y%p����H��s��G���6��Sz&WM�F"0���o|7����=l� T�x��I����4|��ѣ���>� [ͦ�A6�#��q:ֆ�*��}q�f��f#�I{��E��ЀfA�� �\œ.(�E�<QW�8���Y,�L��)"8M؝^��bar��k�����B�ӭT�G_ۅ��h.� ِ9���	�9v�P��V�7��3t;E�<5��6;7��I�=��)?ʠ�v��Π��TN�9�D�Y�`���عn�4�������(�n7%z�!c�S��ݎ{��q����*�	IX�S�W�)1+��U9]~f�1L����u.3j��L�ξ�G���������1S�*A���t&'ٴ�щqV���4�����)�P�x%�:A��{D`�'�O5ZMll� ���.�iЀ�ɑ	���i�p�\�6sfv���N* ��i�r�nxz
H��)ѓ4i��T�%ѡ	x�!Gԋ[��O\�)M%����e�!!���:p9A1W��:�w�C�P2�M�����6]�� K�H���7��j�E�cY������C�"Ć��a�C<�H0��B��h�'Q>���ǯē��j^��(��K`��a,�\8܃0pz>��������7s�����X��<~S�/%[�/��7����_w�:k��ʭ	l�@�ʉ'𘡪9�'�=%���w�dݺr�4z�B��dR��sx._6�j���B��NO���t(��Zhⶺ�� g�4L<E�~#a��w�Ik��'U3��&�ͽR��B�5F�5;M�-�OZ	�{�m��{�`Tv��Q]7-8���	���t��$�0�F|(Ca�\^����z��+�bg0����̌:���<:� ���9=4R���d^g��m�D�r�NrfA���b�eU�4�AK���,����=)�HGH�����|�f���C�4���>��O�������&��*�#��t��<��tZ���h�uΌ����GH4���8��2T�n�b��G#���/�!ę,%���r�B%"�dRW�G�)&^��4����q!8�a��(UU� c����P��J��R������ƛ����F��G7�t�P���
����o��?�J&��!����c��NC��O}�S��~�y����t�ޗ�����O	l0֏'�lv֭;���E�R#�˨�<��]P�����2�-���E��Q{�c-g^:e=����(N�@�ٌh�4���n���Z�QKC��Y�P��.� HDȒx�*�#2�4%��ںJ8�ӑ��U������_���k��"�q��@�t6�w����
�F�����Z'b����^!�u7 h�Q���1}�hJUVOL��4�h@6���H�-C��߳�JB���A���c�<�>�Z(+�3��� �jq?a�D텝�(&�Z&�&��d�p��?�(h�n�_U,2'o���b���ثV�zϭ,6�N�H�3�y�\A׸�"v^Yw�����q	]�Id��=aR:.3�
�s���!���.>������4�b-18�����i�ȏ���L8K�G�K�;�ў�;���7������@�4�)[�N"rH�-��qS�q��7L.����Nk�c�p8s'N|����}4"Ր�岽��>b��c����׾�5H̲e���iD�[�n�O�c��Wo2�HN�(n���) J���>W<c�����bБ�N\�/
�P
��l#��y̑�&<ٜO�I�<X<*Ƅ� �F�q�!}0踔���_,���)���^{���=�q�F|E���X���\ra�Ԥ��^g��c�9�G�w�f��`Z�3�Ȩl�G�_I	%У�4���r�p�Z[����]2=�;󗐡�P
1Mr
���$�eH�3�|�!�d[%��ǡ)UA��Q�r�x7�T�j���y���DU�������H�6�z׮];22"t��<����4lH��S�;��3py|g�S]\ju;�fC�>�)9Q.�!0h8�?!09�f�C7i�	�ӰII1������FF`
o����{��ͥ���090٥N�}�y�A-ٚ�W�;�{/� :�P��ۇ30�jնmۈ|nz�2%>!��Y��9ŕ��o�qn�\_�������M9U	>����Wt�_��ϬY��!z��M�(�M%*xd-p�A���nG55����K��f���H:TR�c?΋�I�U%�\�!�fzB���p"O�ȾK1���(���!f�;K���.���4|�-�l�|eF�ǅEæ@	�͔DIc.y\0Otw��W������1��J?�D�9�qxx�#!��`M)�ϹP�d��F��t)�'����D�;U#�1a�a��QW���F��Ia>��b����L�0"��7���G+�h�p}~~|j
�����fN[ݗ퓄���'��B���b������?�#3GC� n}E<�U�&@����]hR�<M,���Z7�t�;������)��,���W^��{���w�S*�|By��t29e*��|��={��"��jt޺��Ib��R��;n%�e�ړ�*���5��3�Ї~��?��|G��!�e�m�P���y<h�����������)k>22[^�n¸a��������P+����	�f�=q�����=�(����ݰ�����l	J�I�a��,�Z��j�Da�`�l���\q�֠��k08F�P��K���kXg&C�n!e��778/���-�ǃo�ʒ"'L�A]�����s�<�BAK۴i��Ry׮]���Ç��D�*]I�f$�eP�3y"e����gf����٤Ѵ��sٶ�&S���8���`t�x�/�O�H�	z��0�I�G�˟�鍸l)����n�P����tdrY?��&uE���E.[�R<I�JUS�
�)�����kT�͛n�iݺu�5�B1��cG�o�~���.����C���oh*^�:���P��KK�F��n�����t�R�#R�b�k�n�~�5�\��x�ޝ��JXށ�������������Ʉ������@������|�#��;���c�-_�B6E�ݤ�EI@�\�d�U��84P~QF����M��߿W3�w��=�)mJmyܙ��P�(�_}�U\�/�r�e�~�_�|햑��ٓ'��Cz����;�?oӦ7���∻�gPMC"L��b�����K/���KV��=?-�ڵT^��h~�d���?��������K�y&���rR�M�[E?��;%J�/����L���nåP���4I�"�8��8N:�qG)�.�`��(�K�����9�uՊU��}{v=��øӋ.�����F��рkO�1���|x ��o��1k50s(�-R%�%��nꕘP!�������N�!�p���Y\�)�
�������^�(:���w�z�fOG�1Ĵ��(wB�Kr)��
[�8��%�2$]i�['������{��#���g��x@������w����yj�L�0��j�|ަn��ַ��-8�DEi;�-�����w߽g��ãC�Ӫ,�#�-G���Ӵ���7�q�~v�ܹ�0�_JE�'��3�|�;a�����ݻW�&ⓨ���-��f�衇p��������p\a�����?���J�1Շ�L��P���;fX��r�Zh��s8x����ߌ���}���Ҍ�C���~��?�яr�Nc�р��e�tӄ��j;��w�n�W]u�g?�Y�����;��gsd������������
���KW�Z���Gw�RAN��̲���˰�ck�,
1�$Z��ā.�@5X_j��@}>�����������x���p��pK�6<�=-&�c	e]OBD|]�M��J�~|p~~�����xK���S��+CuA�
)�v	=k�h��{b�Ӵ�a/^2���Ʃ�z�!�\�I�6I��":#�!�]7m�&5�4����G���r�Wogb���VI�#1�Z���Mɻ�Y�4ɸ\{�/����O?j��q��'�C\�v��{�7�p� ��(��x��OMN�
8M߾����xH����]�@�/��ϙv��|���R�ޟ߇�-O+��������?����w�����7��F}hh��˭X���ѣ���ռ��˟y�k�����4�������3|���e��/Ji���E����������/La��CRu�FOQ�O��A�V-��'������9q��
''�acj�J�^C���Z��0A��K5�42i��@n��ə��:�f�]��`���B���5+�U"اx�&�*�
�����=�O9|h��g�����M�"�;~�8�.J�k�>�5.Y�f#%� ���\��瞃;D��k�
ؓ��!=4�[�\%T������"�%*POA�@>c	|��tZ��m�e���ͤ����ǿy�K��ެ7p�	��)J�Qu�-��ƍ`�6B�#8���ݢ�(�:ة�@;�������1�`�2�t��$zϷ���\2��8P^�Ԉ�=���Ȩ�,/5�+K��Cg1]H/��	'.nQ��v:Lھ(�fz	M90��Yغ2��w�뮻��ߎ����������Y��g �r�6088:1�/v���+SC{�y뭷^��b�����x��_��W�s'J}{DpN@d���ڞ{�j��6l�h�5�W�P!��jS�������q;pf��g�}V`71������s�e��͛7?��SXĩ�SR��NB����iny$�j��:T�h;�R�'��6�:��L1�>xp�.��R����n��:�����p^XA�Ƃ�EX���p_�=�X�K�|D�����éNgl��3�k�
u�+1�C��k1�7.K�v��^�=:6�ݦ�K�2$��+�s���[G���g��J)���:y���δ�b�jqPs:e/rF1E �'�3��U�"����!b�;"�2�����%�	� Nѩ:w�:l����e<CC�i~؋�� 'L�E���
�~��93�W$%��b:��옚�{f�w&��K�О>��)H�M�۔p��h��X���j¡�C	Y�??���-���7��W��g������;_��Z�A٦��C��N.��f/]��~��_���ӈ�^7�R�裏�%�n�Eg�}��-[�|~�y5y~�����.ܵg_��41�l����/�4�ө#G�lټ�<4�G,o__��|'�d2��1�}�0������W���_�z��?^[".m��}��|�I�Բ(Ē%�Q:�<�R����lk�YI�(s�mO@�Sy�rT��7T�4^|i;$�ʫ������l�CJM��\�=˰LM_�_�]�͢��'?��w�K�/'"�F�`n������w��R^�,8�Ƅ%}�3�JT��p��J�q��zj6ᵝ���իWc���A�	ӣV�U<l��<��㸣s�9�︭�D�\�^q1��������l>T#��b_�̘Ѐ	猟*ǀ���RB��́<Y�29��Vq$��F[<ܜ�����$霦��%水Mâ�]��ܬQKD�I��s"�Yʗ�ɾ���B�6-$N|?�����Xt���LDP�iWV�^V)�M�1H�;�3���l�a�=%dH�hF��D��PÞ��3���Y��$��Kғ���px�7 �������<��7����������������>��_?|饗Μ:���֬]��-�m�w� �{����>����s����i�
y�2̔��+_��k���~���"$�s��1qv�pf��������Ń�v�aq�]��J�^�&g!�R����9����Q��׾����}rl�� 6�|�,Q��!����D�����b�=�{E01X����ɱ�V�:�	�����"5>_y�8���!�ﹰ�bKO��pY%d�_~��M����g>38�O
5�uDR
�b�ƍ��+��cQ����3�P�+t$���*�J������/��\��%b�B!�.B#&�4���Y�2�5�����d��~�	�'vF��`gf���V|�L�:[9�pc��sZ9�Q��
���@`ޣ�?��(��aU���-���L�K̮h=��ZkP�K:%����s���F�{&p���ٓ ���Y��%#{c<09�#_���)��z	�r�3�@��`�����[	)#��É�O�UC�������d%DW��O���3�qI��/[v�����_����q�7��g>#u����Q�� 38��
�hv��:G[
\"(�.� �r��z*�7�tD����P.�RV����Vm)T�|ڪ,:��R���:M�ٙ�|�o���R�`��1�����U���c���%O����K��^z9��Ϟ����?�o?��U�Wb��=��/m/��}T���)���a!B�.CJswh>VHP�r��}O��O#h������������ a��F���#��n��n�V]6XȨʸm�����U�6�/T�N��f�q���_֟���K��4k��¾:��x��O~��~�o���#�(J%'԰�;oַ�f������ժ�+V�'gO��-o��tcn^����<��+*Ž�L�����T�����=l�k���2���Ri�B�Y�a��.�/�Mʹ"�'�t&�Gs��`D!�ͥt����5�y��1��S�K*�nuڵv�ʦ]�ZI��5ɰ8Zԅ9X�S[m�"I�o:C�"���a�;~K3��C@+C+q}+��wl�!���G秔���n���mU��X���#�ՠ1�k���f��CC<�P<�C
��r��pu��&L��P�!���)AK�Z�����q�)�o����
��r����9M�i��~l���
��z������l���
�\)��V���)ab��6;����G�v����Ç���ꫯٲ
]3��g�ulnn�VWs��l�//_�~~Ǒ-[�ÿ�:΀��/�VL�M�	S�0p�2��M\^�J�Ga��W�W�g�A��+���s��t�SS�\�/���r�ww�ر���-�����JTG>KU�3F.ǴS�#63=�Ӆ�t�h Y?y����Rt[Ra7�0�gh��}��!��P|���`���΀R�τ�,�V���b'�v:�eU-���v�aT�2%��;Ђ�ɉ�+�qe�#C�'&p�k�Frـ��Ҋ�j��H�LK@gd܂��F�l�8�)��/!nĬ0��Q�)�9Y&�z�"�J\�N�����FЈ;�,F�J�l�^��W;��8������GN`����0��EA&k�]��P�=8h��w$r�x�5�؝�����m�E=��6�K�`��MBH�{�.���V�MZ��+�뺺0�Q����
7s�uHP��rƘ�:�*J���)�u�������@���/|�ﻗ����U�:ׯ_�G\^ZĖ�X�Z�o T�����^��x�̢�0�����=��(K\�
�u0�x����VnM/�ŃA Ṋ�L!߷}�v'\�^85
0ހ֛t�N�8v������Avy�R,����k�n�1�WFR����׿�U��w|�'�99`ܖ.Yw�8el�>�,��ˤ��l.�ɖ��EC�'�M;r`bYI��}�f��t ���B^?rxO�� ����1mʻ�J�)��}�|*�4�_y�ɢ914�����t����A�����3��ϭ(
wj(j�;�E�BBc�Q�o9��b��i!�6��^��8����3,b+P� .Ζͅ{�������2�:,-B��sCHJ�����13��&�Hݐ�*y�&g�$�:N/"8D)W"���xB5v�}�{�W\E���#nL��?�+� 1y*Jn����&,J�
%c��	�=�^I�2U�r�ժS����IiD�|��ז�D��mI�C�9��(��-�w�w��∎RJp5��\Y�\p���N�����<��s�B��h���s#��r�$�ڶ����u�8
�Pepdx���v�6<6��&^zdZ��f]������C=��c�3ӹ�Ⴧ�?040X[�@y-��!>4V���K-�P_<�jj��|�JYf���B#��'[4.[I��csa^������w�E�K���,�5���?L�Sb\ԩU�G4<6����Ǐ�@t`�X��ٺu+���s�%R��m"���$�����u�%��駟&�]�p��p$��������y����UQm�zxxBb�g�,��,EMYķԢY��Ӂ��!j�5h�ǣ�Ȉ@[I���-�:ujdx�,[@�18rl��=��a�Ej��Y"
�]
�#�RÒ�q��u"�	5�B@l���CB&�I�:Cm��@9��S����q�9c-Ӹ���m�� i�'�L�ɨNb���"PV���j*w-hĭ��i��t���?����~6�r�����t.�:;;��O|�O�iH��T�*u�\��y\U]��A9�L���L��3�� �
U��!U5���x������F�ֆbD������?_b{H [
eBI`�!D>���)��S���c����/)�w��
[���/<��"�8�ǎC\����{���7Z&��*Ҕ�T����`ȿ1004=}�������v���w?���\z�ʕ+V�زe�ƽ��|N������o�Tfdlo���e�>{��k�����#��[��я~��Wr����	1�yŜ��iRjfm�A躪!�W�����C	�N��IۦYz86Z2t8��N�d�[���a�x୘,i)#�Qjծ�TE�����b̀It�@�W��v���G�ٹ�Y�*�y�637c��6�g�����������A����]��n�Ͷ�/��*U��dөv��q�ju����7�1q�O�:��,[�Ã�/`'�e�x�K�F�Y�Zn���z}ڦ��f��X?���ӝ��5�Yj��&	z����u�T��ntb�O�B�P��#�
�N��	ȇ���F̉W��?ʚd�y<�j����F)-�Qd=�%�#��R���/�ZB��/���e1��&�?���f.8#v���'��4e)=��8җ���h��������:�G#���4�sL��X1E(� �F�Z�|�L:��gp .�x��S�_|E��劘z�=�q�b^�]g�ƍ7^����֟�
���=>1sJ!��!���_<x�7LM�o<����r�Z9��C{��q��؀��ٳn�z��v��;}�H��,�,FJ�ꄒ�e��s�=��G���.���Ss�҆U�X�\�\"�ů}�kؑM�6A�@�Q�aiidl�c����w}������~����|�Q�;��~Bx8ғV bL�.���F��=%�L�I�,�A�~p��4E�,�L����U�T�/G�-�S\��ܒ
׈�d�Ԉ���X�C�3gQ�4�Z�������V�t��������D�R�e@����J,]�b�qj��w�N�d:M��ϥ)y�����G��J�m��d*�`W�zD4��k�U&-�m	 @���"w�G\���qC���骚��ġ��=O<��_<��f�W�<ڠqT0K�O+����y���ӕ�.����|ĳ��ಓ'N\w�����ĄPsXL��\��RVC �������zk�^��M΃I��Oу밼QX�֤�zU�~H��a���A7�>;%�_�� "ݱ2�{�}C��B0\}�����X[>�
��!�u,�U�\}��w�u�0'o3$�xG���@;���;|�F�m�x��͛q�p�����OM��H,[=��,��w�8� J�mƩ�Z�Pj#�\�z���G~�庭0���6>>�eU*5Bj�}���ԧ>5�l����6���iCG��w�����������Ї��#�0��?�q���HW�����*�<=2>�� /!�f�\��(*`,�/�u;MK�Zi���Ù���m�]U��r��64�A������&��Fv<[�J+t+���0�Hug���u�ۆWIY��k�E8n���R�Tx�tv�������������l{�XO���)9��4�+���P�F�|�h�b��r���{�����V&�׍xh�ۘg��L������n�������-��f�-$��$�j��*�2��+������E�֬Y���$���1�&�^S�0�V�@�D#�m�*���C:K�!��;�isێs!\�����n�%)B���l�m�ROot�&1�,	�t��Ơ(��;����<������u���������~�����d֜2�U"F����\D�enn�����)��:�4jq�T� ���u��=(�������oT��ʑ��淾ipdTg�<ѱ��n��T^|~�3䈞{��?��G}�o8k%ٰ�����U�۞}e��4�z��H������p38���{����?�Al%6zbb�- ��p�O��_���a-��x�K/�$*9dn�l,��h@1���җ���?��}�{��?�q�Ӷb�u�	+�����s����ԁC+z�Y%!W�CX�i��9gM
궡�<A�Q���T�QuC��_X�8b��"��KO��fa��pȐ[2�QA4�&���7]�1dVKm۶m~�0�8�X0�޿T]�$�޽{���g�yfhh���~ꩧ~��0�Üds=����v(���b�T_�
�S�R�����U8�8-k��9k�[�����Q�)��CE;y�������C��:5-���]yGw��qj�.���N�2�<��*D���!�X�?��?�����E*�gvC���O�]%�����*�Y%�cb�S�Yˌ�Aޒ�d8p��mO<���v������|A�r�2�p����W&�GM��d��F"ZL�3�'�	�`e2?�����Z�f�7��S'N ���O.��o�!��L��g�zl�\Sx�8G�Ї`�Z�=����"��z��<;"х#��'B�0�>�[�..��]�Z�Q��|�G�}�ٱ����^,W\�X����m��7�Є}Xn|ǟ~����/�4^z�+WNMOn6��<�T�AD*tq�}���ž(�%�߳�檌�t������ȅ;�*q%�X�S,T�V8��h8KX�4��rp���b�D@�~�I�m
�a�u?՜�"4�;��WU��6�8h��Z���.��B���K_�b
�Sz����j3�f�vY)�EJ�Z�C���3�����x{�ŗ�O��4�
dr��4WD%�V�-.+�aq�� p�|Ǖ��\+���.�*�0l0p@���Eui�F�����嗶#��l��9�5Cw:�z{��E\�<?o� (�a�0�on�k�V���ur�#h�гS䋲���}"����C����SB>��h� ��0�T+��l��8���m�t���n� /#m[�ͺ���U+u6P��2\Tw��OΈI��!4��j�w�9RJ�\���瞟�q�0�+W�M;1W�z��}����L�-4o3M��V����=?�	"�u�V�I"gDiLO�ر�U����9P^
��>˰��Ů���4Vԏ�t����sز������m7,ŽB>�aÆRq@ҧx%W(
�"{Z�~�Me��yϻ�50<������+�H�B@����10�� �˟���OI�<�1%A[D�+0e=<T�C��X����d��r�����g�3&EH�k�����`���X�g	))�P�X����h�/~tt W�뇏��	u����^躔�~0Ӣ���5k����7.M7s��zwڮ����;�1�rWE��QLM�%.���$
%T�ْv�*KvQ�'F��)��1[�z5������
@j\�,X^�,��'���PB��Ek��K\d���˗MiI�9��+���S.6P�-���:s~�B2)�p�A��33�hYgr��;w�T�D���"�<24�����G/���H��l0}�O5$���P���e�Dܝ(% ��x>3`�r�������څ���[�g'�I5�,M����\<xp�֭+V�T�ڵ�WvMOOw��5k�t��@��(�Bu=@)�j�*:�'�ﴝɱI(-���6&�Ac1�%y5��vݘāN�O�%�0���1�:p{�ҚYPu&-N4Sk
yv�
]I-�����W�׫m�[�/醕�+������M��tm�T=�\+S�Z�YL��CbIM-_�?"�;%���d�T*P�A��찯�]���#�t"�`<@�g����ӆL�\��4R���u&��3ʄn��у���=y�ٶ�`�F�^oJyD���Y+EӬ4�(��[��/�-.V��ƽ;>S�7�>8����\�qD�>D5d��ە�Sn�c2�D�b*K�°$ēNH:�I�G;=FZ�N������k���`?N��={����C{�P-�I�\��I��ǎ���΀�����o�ejr�����l�,f�v�^",�Z'��$ÄK�6Cĕ�G�S ς�*�tG)��g�e%�1G3c�@֧�~���v�{ᦋW�^7��p�<�I��-
�G��������q���I='�|A�	QM��{p�"�U����߹���C�Z�ܲ���P.�hsw�6�5�ՙ�X&��H�o�^�(��T��˃�gt����U�BS�"7�Leb7M������z��2KC��o&#&�����L'��V�\xᅈ��֍n5�`VJO1�2�r�\9�P"]t�aG�Q�5r�ͨN�\Y�W ��j��v[���Vqb������YZ����/�����Ple��)�&�U�uX��x۷���o��Roa�4n�L)о"�o��y��6-�:�+5�e�p�4��5k���zL�/��^�F��"��[S�.Ī����mpқ!��v$x�*���5�V����6m�Ԩ���~��OF ">�B�ݻw'��>i�M�)�����\)튐Y� ��M�k���-�V2���Q��
f��jn2��%i4%�'B#�
��T���E��ױ`��	X��TY>-C}k��UBk�HQ���֘��ѹ�#%�44D=��t.�L|���ʭȭ�,2ġ�"�bސ�����4��K)&�P��i�d�tV�ɐ�I(6[�у3k��}G�V�Ŝ�|����A�)w���o�2
B��nZ1읡D�60 ��B�5�b��Q���b_�XQ��H}�"C��c*�)���Ѩ7��L6�[�#�g�߸z��s�o�5�T�q�D�Z����������ae�%\����e�`��!B���N*2�R%�"���:2�	��uk��� <��(����S� �a���-U�SO�8ި�<G�f��z�,�_��M(����|(�����hZYZ���[��B���R1�����a�fN���ٕ��t�t�T�=����W{�I��w%	.�p��̾�⋫V���X1I�V��NQ���C���2�r}�vG�lI���YOg�H�0�Z�R�DU�+�
ek�P
 P�Ͳ~č����e�옠_�r:<1D�TĬЇ7d
��޽��1׮]��C�)�Y��01619>��5����,ҲC"����8��c��G�i1�e7�|��sIs1��D��� T�ԉ8S�Ձ_344�n�-�d/���?*/�;Y�D!4hJe�q���Vخvj��l`�q+#t�8ʄ��Ʉ���g�u��%��+��H8I!~��XV���rX6Q�t��R����������ɀ;��d8B������]>��->묳� 4����~;5�R�Ѥ�����N�O,[6zpId�)�E�*�xf��sLLL�|��+3D�!|��)x��@E/��wD���wȍTX0\��}�����qnܸ��ѣ�qS�6��(.�dW9�*@h`K��)���a/�KiO��&z��Q���Z�X�?�{)j��|�NDI���l��M�mk���(BkH�^t.��@F���;}�Cv;�v�R2Q�)��= �]eN΀�� �T�b��%�D'�2%2������6�?b�Y���*twX���co���3Ϝ8A��UW]E�A;�����o�����4]�[��˃�>p�03ޙ���g�K
f12���6�g$�'��;<"�?�#����@�x��_P�S`F<�)�!N�$�z�U��B���JL;���-�]7z8�o��B�&�<8�*�n�ɳ'8���d�պ�z2h2�)�∜t�j��a�AA�8V9��𘡹�������AX���H��f�ڔ���702�Nk�Zc�����	�%���|Äs���#&���Lr���:����c���C���l�a�98j�Y�N���Z*?ҐU(���t|�ʕ��L��z充R���ކ
����<m&'"��):����؄��*,\.b`�!�=LD{�	 ��h2zS��)�!M����$�2�PR5�>�PC�Za\��$�S�BBL%>'�(nlu��v��i6�C�SMy�ZdS�{����Ƿ����� !���/�0��������Uƅ�G�8!D��>��#���	d�I�F��T�����٭�^��O���肋��كF�dlb�0��Э�h��MAn��\d�x�j(�Հ��7ƋX���"%�#�"�2+���vB��%�gV�L&+i$�����i�A��/��'�-���Ӟ�h� �7���E�}FCҬ�~�����'��kܪ���D��%�I�I3L6�I+7o�J�R���8��	�jr=�#-����A�:g���W�;D$��J�
�ǻ��
�.�m�Q���©gW�n�!_Wǿ?)R+T xlb��*��F��V���V��	۶m#��,��A+�a*��Cċ��m�ry��;4��T"�帗;����bJ�D4�äHIt~��B��;B���n2s��d����)��&2C2�qs*�!e��Aq���/�w<y@��W�_w��b`-�K�Ԅf_u�- M}25U��⣚�@g�]�k0�F��S��@�g9��((1�s�Z�	�,�	�kR�;��P"�o`�yUS;w�|�{޳u�V�~��^����<���ێk���%�u�6(�ǳ�K�D��	�jL�>��O/+A�7�I��U!H��v|�@r4RHNJ͑ؽ���J������|�Q�pJ�Ռ�E\�$���լedRv��T��Y�j��|ڢ�JM̈́��7�fڢf�v m�n6m��������HP7���nz��#&��j�6���JU�F��Fpl����wc��Cr�i�l��	�
Ť)Us�5"��pl]ݴ��٥�_�50> ��vyԮZ]�.�g�;6S5��睰´S�idp,�Z����r2�ce2#aN�:\X��5�P���f�5r�ɳ���}*cg�nC�ۆ��z핗�w�d����RC�Z7-߰20�j6BM��L��% �Ҝ����v��4�vM!�mg�
#���ZK��L�H�-R"x n�9���"�d9^J�$�'��a�8��3i�Ne�d�v���U���ȉB��[��5�p�<��D�L�p�[������w�}�T��zJ�W��@�rT~*�=���CCA��Q�C����$Dx72]�TEǆ!FS�*b/7��V_J��]��)�ȏ�b���D�ڮۺu͚5v:E��M�� �l����=SkU+���[��ڭ����|��X���-6�So}�['�h���6�8��̜�8|p ���h�ԯF
������Ӂy�ЮK���R�4�J7��ˈJ��<�C�s8B�N]e�:cg��t�Fy��b�m��^1�;?{dp�p�%�?���F�2|[	R��!Gcz�I�������f� ˋ°���<*(�38L�>�i�4��>y�L��I����U��pO�1.���
�+�ڐf	�iA����1�H��U�@#-x�Eq�Տ?.�م2�=��˗?x����Y�x��.Ċ�G�1Э��!���y�C� �NW1Om>�s�/�L��_��A�-<�n00==����K3<t3%s�p���=�<���-b�/|��M�Ҍ�W�(G+.����#g�fCh�hx��5b`t��a�H�����~O�����De�p���^����\�A>�	�dI�O1T�\ɚ�	���]�٘��jm�1m1���d�[
g�x�K_����d�4�ok:��Ѫ7�;���?��6�9N���?���
eq8�}����H�����m���?���b~n��/ҩ@Xv��gO.[	��u[W\q������M��B)̤�98��C[,�wC�Ik���]7�,����@L ��2`1���`�a'ݷo��,d9OKs��0h9]�2�n;M�@kr����0�YG�r���)��5�9!���F�����J�����g�T�C8��5���n����쫑x�r��tV Yws���BK��&������r�Ru�ֆ;Q�k444 ;s���K���=�l�t�ٔ����y�S*�Zk�2�#�`Z������9w���d�Z�J@F���pc�|�I�7G��|6O�GRc����Dߘ"w���ǨE}���� ���h���ј �1��@̞Px�ϲL�kehl�9�$����������R`�u�\� 밡&?�C��1�5ղb����{A�+�kJ�>(Y%^�	b^v>����dIB'%<���
�*��Z���Q���r
3y���'^ij0"<.H�ǥ�������mO�y�G�fR����q�C���+(���x�	�����A�ޠ��������3Gg�z�$ǷW�\y��~�_.\p�?��؅��c�zubl=WT�4Gf��� $��ݣ�O���C��KKT-��1�RbZl-�2���i�l*����p��Qf������p��t
��
�d�2#�Iw�jQTQԱT]��W/c��,L!�12-��-z��C�֪�GDA�|E/6yX��2�V��ǣ�|�¨'�KU��I��q<�ז%���5�\C��2G3�ڴw�=��.��2�������<`����`�	3�D�b�n�,ޏח����S���<1B�824�cǎ����u��?Q��6�M��C��p�������n·T��)�J�L�l�x�%e�0:�A�u��.	�H~��aj�A"e3��ٍP��D� ��`pC��6D��'T����]��[Zp�A�A�oT�ʙ�K�+a�'=j/GN�Q�y���-"�%%0&I��#�i(�$St���
w���X~��?�T����׿�������eS�}�e�$�V�Z�����`d�oߎgtt�����Ga��xR� ~b���5Gs�4�޽����,�}�3�䀝�ް���'DN�
c�^�|��.��$�y(��~�|�I� ���1���T�IK-���)��&��P�N���+s�|�^'%�*DY_�_���w�{�y��W_����m�C(�l+8g��h�x�"=�M�k�P�3�@�&��2b���*�J<�]�(S�x�8K��Z"8�<�[f�1��x\��mڴ)�M�k�%�z��o� �����l�44��>��tZ�342��Q���U6>�����ŗ\جU�#�lz�4��A���c�C�s�b�l6CO�z�t�ԩ9M������O�qB�=�\|9#��95�y�#��T
#H$n���T����9|l߽��O����H���˩۽�۶�vˇ���nf4	$`2�@�4���Fʹ��daӗ1�^>�P�P�e�ĉVl:�4r7��*��8��d�|� ��X⟄�p��\�	�@$ߣ���ryM�lD̈t�����C
1t�׃��IJ�A���G�)k��UR��6sbr�57w�E���)�QC��l�2��=�(�-���ߝ\6�����O]��(�Ν}�ys��8�k�=�8;ߗ"3�(��\O�P�aL�m$u�>������C�^�H�Rہ&���+�5�����0M@ 0Sull(����HY;&����Jy)��4̓�N����{�'�At���[n���]h������o~�[�5����|�+�>��%�^e�Ķ�͂���f{��lj�!T�@�.���mO>%�29��/�;:���s��<�Sc�ӄ?+�_�� 9I�R�_}��W_AHE;w�4������������#�wQ�#!2��׮]+�h��|?��_?�݄��g[�:)4�'��9U����\�i4��C^z�%D��^~Ŧ�7X�0�Xd�E��0���g���.N��%z�|[��"U7�(�wZ,��niΙ��t�cH�Yqo[<�T������ӧ�g?4RO7�H2<9��X<���JBs&yl�	��d���~^�Ȝ(	UJ�*ܼ��B.Q�	y&1$��^~�e��C!/�{��A�?��F� �z\�ℹ�}�#?���)fJ�b�Od��僭&5�u�dY����t�.@��a6�7�t߂�U^�j�s����;v�mFE�b#tu>g�	_](���^r�&ޫ;^D�Z�_���Y��q����c}�CA${:6:
U��p���uk7|��ظ����W_�w�R��Ͼ`�R^x�-��ᦛn���?��x�g��[��xp�
M�뮻��?�я~����謍ݮ�k^q�e��_?�p�m�--�q ꔗ��!+Q�0��	ܞ]�^]�籕\�D����o�h�7nxlT
Ǜ7o>yr�駟�?��^�|e����C��2T<�p�����h�/n�����U� U�z��?y�yj&�ukqe��K.A t��a�;?��##C��8�T�X�bŦ�/��k/mߎc��0?y}��C���g�{�N��3F�w�UW]��,�kK��R]Z8p`�
12A�}�aZvJ�®�/6���!��'�sԘ=�e�O,��Ux�'f�-H�Mf�^�HO(=���������*q�_�i���s�����ފyuq+�U�s�4�V�>� ���z0��*m��ʱs��<CRD�"]teE@v	��kZ���(+��H�@&�<��3=���r�U���sNU��}����TWݺ����sޓ�C���FF5�L�a8�X���S\������PRW�S�+�XѶ�f������55Q��#�<И�BZQ��P�Bk�$wlCѨ�����0x��9�K�_0�ǅ�U�!� B���o��ƛo���;�ؾk�a�+k�̙�V�O�E�j���?���N�5�H<A7��S촩�������q��gΚ���DB�;�y����SO=��[�����y�4nC'�;z�H����p�?��Op`U��!Ѓ��f"+.���C�����C%5
<-4��y�P�s��yu�o�޽n�!�k�.l����|� ڜ<�T�|�SW�d�r�.�Sᚚ�~�4���+a�'��(/�rmܰ����b��c{}x3���O?ME�^o z���q�!�q�[tN��+%��.
S��z���_��V=vt<6����҉����^޻{�be���@Ŝ�x�ytl�����2~�'���Wj�*� ���Ь4뻯oƌX���o���`8��K/m��f�M�<�d��+K��V*{�,��(�GLY��Mw�(O�>)&5o���S����@V3�U#,�Rl �E�@�ǆ����WW�q��=s�6�ZV��F:��; �U�ƴ��ԉ*�V�y��K�Ē�9K,ߎ���� �>HͲl�垽��։�B
ʩ����������n��DI��E�P1'�Ǡ��%KN����Ł�9s��}��}������N_u:��w�a�.U��C@C����K�o޼y���=S{ҍٛn��p��~�m!)W��\����q�_�Q��-_�q�8"'�7nX?24LCB
�S�u�yk�
{�|������m|�Ё�-�fy۩	G 0>.C��E͜5��.��f��إ�y�7���#ʀq�A�v�1rEq79�I�Mv���Nhzr���Y[������d�m�ݶu�f�57��E�8�.L��ӏ�:������?~}���Zۺ���g
v�/^	a���`ߠbp�4γ��@�EK<^���KqW#��W_[�W$R#Sg�8vp����8� 76B�U�̇�C]p��p2��W�Z!}Ҹm���w�� no޼�������K�����ܾc��m]�YK�Ђ�W�e��2��ۣyM��i,����ῨB�j�+M"�p�|�O��Oe��Ly?ty9�T�P-�i����J�8��Rx��p#�b�����N��ܔJeثTҩl.+dBx����Ţ�n�u�X�x�آ�|n��)����+��d�37���_�hW���tM�"z1�	I��0��0�,�)�&����p�H�NS�L���H<���$�^����ܝu��4T����9�q��_h���}~��_�җ�}�Y�
����)9��U�.��
�ޭ;��y�|�M�rkS��ށ���݋�-V��rt����>�l���/�,�-���$����~��3�c��w�۶m�#���[�bc(.j1)�_��,^�`ނ�&-��2���5��~٥�I����p^��	<�+_�K�\4S�:�7#�`������ڛo��H�H1C� ��'b�@���[o��H��ڹ�?�A���T���(p�e�]}��.Õ��
�#�Y���̙E�%)�GGp�X�i�fe��Z��R�+�A:Tn��2��cw�����V��P=�������O�T����zzz��:Pͤ���C�?���I?�`� �Q,9|N��k���I#�	�;8B=�D�2�Yr�^w�*��^��HPM���4�琳�+�j(�3R� �x��R��:2�ExJ�ʭs�DBF���[%�WT
��S[$G�.Nd�--2�Q�\-����>�R^�������w�_&;��V4�p/��#q�jpK����}����f���7�����_u��{�D�a���cP_�ۅ��9s&4�'wG{�0��$��W��={�w�Fv�ԩ]t����1c�b��X����X>���I:t�hDH��e˩�Э����j�p�����GM'I;��>hn,�|!o>���#G���i���@^D�}�
���6(!� ��ci.�m�-K�q�L�p�ɼ���6\z� ��ń�)�Ի`�i��;_{�|�a�J�000D	��c�r$]S{t׉{�w,��� �0Vx�h��`��^<>�#�{lt������7ַ��Ju1�إX"^R��,���@b�A�{iR@Dlr�{
o"�N��%ER��)����(2���7�H���8!a��m�Z`�����D�+��OT��Ŧ0�0U$<g���.�XQWg��4e[���T�J�o8͔�*WZ����4�\qb2��	#L�8��qt���PŹM�!�&U���`��2�v���\���Z0 U�h�C,�&՜夈�Tꢊ�X����Fh�T]]#R�X�T2�7#F���Kp������eDJ��w�O�����J����YBu�5��ټ�����:�AhP���w��﬿����/�m���ű��)��lB�p�1�W�P����
_r�%����^���ށ�#t�a��YS;:�7}��0�>0�@j��R�.�����+�\$b���+���$$�Ax�5=Q�E�(ν�3�<��;�$2:�Д/��P׆����!?���m�Å��bQ�Iw�P��������~�S��T�.
﫯�8�P�HVT�N�<)�� �{[0wd	�(�f���/A�8�D�Qw�y��w}[�
7�*��N�s0J&&�͗�8׏''��@I	?�w�L�)��bH��nq��3W�Q �E�	��.�r��4gȄ;�����4.���#�-	���K���<5IE�s*��4��́|�]�R���V�T�1��P?1#ުDc%<+@F�Q��w�^���@�Q.�U��֪i�[r��T�6�
;��U�0&S�@�S�	N,��)���J/�n�x�,��4��Ϥ�\�x..=�{�������_8�QT�IGJ�U.jW�����c�]�si��@��t��xjؒ�_~Yz&�28�-m���~:��Ν;! >�Y�l�O�t�R��=[��.S`�iӦ)ʛ�D�m�S��4UƳ"�QO�����c��ٳg����y��9��<�?�����P_�{����&�.SCC���_��7��ַpm�����H4&��l�3�c�Cþ e{�x3��\���A��&GD����;N����?��Il�M� yZ�n�il��B0����ű��o���d+������ޝ�v��Eﾳ�����V�X.*�q	��kՊp�w��	�o�����fG�!^������(\V,�5�T:�а���R?���s����U!�.�@���d�}<HI��Jm
+%UW<.���g�.��ZA]sJy�W9I�?�Jr;�[Nв�ш5.�;2��IcՊ�(�XjS�
��LX�\���:�#�tD:����}� �\@n1{�j�^�;�'֪L*���.LCC#�\����0�I_ 7	f�4h@���L�ع�kxg͚#�	�Ã8[N{��y�h�I�S)�H[{K(8��s5E���E�h)�m���tȗ�#�K��tb�nkk9z`綾}�7}�\_� �\
@���pm�m�u����7I�L�|l��E�!jy"��MUq����p����F �)�N (��cW��#��5��6P.:+�q��<�[x���Ӆ똸�W@��
��/��w��~�G�gÆ���Ӈ�9s:�K!�O�� QI(�.�u����syb��uH8$�Gy������o�;�=#>V�U�Og�i�ౄ&<ęx�
E�X$Rs��A��nٻ�P�ƚ5�������g]m4��f��� ?6_`~k�~�7/��:���b;q�)Ŗ��?���K�	B�.�zI�AJed�U�
j񘇪�5�̫�PqK���4�	I�Kܒ#.dR<�r�X�&�O��k�Տ��^�,R�L��JPud-yr��Z��w������.y�(�2�L���`�twoݺM��j�Ͷ��a'3��ո.}��r�J��}�{{��mmk ,A{/s���b97���'-J�+VO�yM���F�rI3�+��ԍ-p����\�v-{���Ç�
���������=s�|��_��g9��E�0�,�TJS�%Me����}����8��[<AI;v�=��:Ӛ9����Pb��zMs�5��M�G�7�����?ًK<��s������_���?�r��T*��x�bi��-x�)]S)��������D�C��%���Z���n��w����O�QkjC�",Ǒ��?Yw�I�n��bQ����g��o��PW���߶c�v�ϝ��Z[F��cc�Dx�A�v�ً�$&>�'�q2s�dl2�3mک������M�ڳk���˗wv��2y) O�c�4ZCU,��k)�s��ԗ���?���A�W�E�ѱ2'�W[$��&	\�+�Jk�:�0#:������YS�2�+�L����T�41:f���+7�daLy�P� t0�#y��C��6�[aj\��GC�Y��e�"lr��k\k.AA�U	�:�"QR1#�Q�6Y�2gz��u�T��}��M�)����XT�b�XB��q]1ū���p�:�i��d�n:$T����S��2��s!�Kb�{�<ߛRP��URAq���5�;�I=zƠ��~���K�'�~Ό��sN�2a��hk�<C�jB5q�ד'���o�u__����-,fX�Z;�̳���P��MNƉ(���F�Ѻ�:��>����1czRIO����:(Џ���Gu�w�r�/i2guH�D�j����'&&/����ZnM$ĥtP7c�MMO=�ǳ�>����o�b8�T�J2�)Ox��sլ��O&��������͛��n�K���/_�b��vX�G��SP+m:=k�,���w��`�G�_~9T�������6y犥�?���A pK����ЩA!��'nr%-Ⱦ��H�w�>�bŊ�8��(r8��������pz��
��l۶�Y�3lI��X��秈�#��)��&<˛�ކC�;��tiPT�Ds$��!�#�8��4$�@�J�����L<eS���~�+w��}3)��z Io���ڽO�T=��(��(�L��R��NM�$6طT�)"á�Du�����p������F ���'���FΈAݛP���w%(��f�Gq0�&�N��9s��Y��ݶ��H����]]2p%�#�Q"g�)����s�/��Pu���Ԥ�(X)�� y`Λn�	(�~��$Eq��1��$Ӌ��=�һ���[n��?�o���5��d8���}a
D�¯١�OuJ'�{�����|����p��� %RK�.��k���Ñp ��TߩW׾6g����q�p�UԔ`4�;�u-�P��׾�u���ﾛo���_�xr{j�2o�M�N� 	?u<���E�I�x��e��y�f�+{�w���.���}����%�H��7wÚ�5����~ΒYW�t�}���/��1������s��{��S**����6��ڛn9y�pѢ,�agF,E8mÃ��=�k��0Qf�LY��?�e�����U3��q�w��%d�a��:%�o��C�=�/�)i6<�ں:�?��<�����a��;�<l|2��^�x>vn�{�->�B�.:|�T(y�^>:w�Є	�7�S�u!���Uy�߳� �+%;O;\���Ѧ�(�U��'MF1��T$C��!a��Ё}��Zu7��/�2+��0.S�5P\m�ih���S^�SC�=˪^�z��W��z�v����p8dRy��T=�bڶR�c�DL?	C��(NZ�J����?Ҭ���}��_�`Ӗ����������LE>Ǔ��5�	z�����Xq���X��?�:7Զ���?���p�����c���$�F��|��V����C@��a�Z�Q�F�.%&��_~�E^Qlim ��0xl�2�?�$:N��tu:v�*dR�����i:�^_��3/��x��%�?1�8�����)EW2��Σ�DQQ��X|��w�̛�hѢ�˗o�X��p�B	'ǌ#��v�y��a3g�,�4�%O@\���וg�	� ͍/���>�~�������8`�/�ַ��#e�YE�P��-��U���w��~ٲep
h�:G�!� r�ebl����`�Νug�b2섴�����A�$��j4n��z�Z�A�g�?���]��8
8QR�ЭP$M?������!\
y�e�=��ol�n��3ɡ���,6S::.��|���H���mdtZP?J��y�����̘1ϸk���������z��|������K�T�ޖ*J�����<�x8��}�Z�X��>�*yR�
�Mi��XK,�T-J�VЬ�ز�S����w�f�U���6�-�W�)�uE���%ԃϡ���NW�I-q��A��Ф&&.��B��x���ϙeيW���]�֍Y�gc��<��@0L�1�bk�L�'&xp���+x�V��.{����{�i�Y���� �*�QI{�v�p����\s9Q&ky<&Pt<���t&��(�ɐ0nBg�=�Y%{�J�Bp��ӻ�(":3�ݠl�֭��@�|�h:���*��n3�Ǳ;���C�~����Q�8�@�ni%ͥ�G�p4o���7�xc�򕊪'�L�����y�ah���Sw�}����ϝ���w8W=��8sMw�x,�&j�B����̙B�A$�����D��E���LO���H�4��F0��'S0��p~�sk��GJ�r�i��{o��q��9�`~%];9x
��sι��oв�G(:�a]����d~����#�p�rNP�
�y�c�"��/^�З�X��RF"u�lM��J�^��k��y�����q����������1>2��/b��M�i�I��29���G R�Zfa�A)��g���*mbє����8j)�y	k��p��B�� ��(�T�.�C���9?){������@� �-19NW����ke��2���A^�$�A̎m�D]�Q�f�ĉ�T<�=����褛�@��h/�,�6Ο;��/h���3Ͼ�fm*C�V�x�6].��B�I�14|�����\:[z ��Y����hِQUW$<�1e����DWk�XՍ7>������<�}�cV�j�������+W�\��ۂ��7�nڴ����dA�ܜ9s��a-���%��L��߿��ᱝ�ƇN�|��H��p��]�W�P�K�}�c�h��+��@�*���(����5�<x��3V�������I��s)�P�
s�CCc��A,���5�U�&И�JЎ��J��-'��'�*@�E�r&���wf���:������9<�� ���.��R�&@�6Wm8pw�+oI6R�Wv��g����^*�5�t�ͬ�!�ЋX((0��Z*W ~�,�Ơl��@)5�G�����S�,�X�q��*�=���}��ёq�6��+��P�8���a�&s����J����>/�d����fFŚSN�2�^&�@J�H�o�bF��r~�OJ�D��V�����D���җ(�0�`@�	qf�g��.��*4vgr|H��X�W�����+|������MQbrF�T� <묳|��=4$T ���� �0���C�&���t�G�x
���t�N��I�6�C�����c;B�c1]�	 R�a��n۳p�\(Ǐ6m"��˚:���w�M�-���W�<���q�9\� T�(gi4�2�u��lf��*	m!q55�P���E�i���t*�p��=���6tO�>℥ă��;v�8�{Ok[��/�Db!����a��E)���-���<���?���~w�-7.[�b߾a�	�lW "�4IK����rӭS�9�`'�b��������.3?:�Өv�DoG{�d���`��D!�8UuGG��X��w�����Ǳ����;@�w��2�%'��JJ��鷋V*����3�<3z��B0(�lk.<�K���(�8�XN�)*q�|�i�z������}�cS�>
$����KE?*L����n���������y�C�D��18��D�C�4\$YTΪ����m˱�1S
>u���M1_� ��1U�J�;����T������Z6W,u��Y�E��qi���<t�S�j�YQ�U�OR%�ɡ�#��%u���P�JAx �R�]��Z)+g���a���z��_������p�_����9����3��Ԯ)��5�">�q��}.ob"n���#EE�f'+F�D6�P�>���iӦ�}����dg'�3M���39W����~e��J��4�S��M�>�Yg9�����:t�_���|p��%�v�hh�"���w�yn>,��ԩ!�G����`ά�3��c[�l���3��P޾����`l͚5�Ɇd:u�CQ�i�tIj�M��U������gir �C\�t)$W�ˈY�a=X�_� ���y`�L%$40�l�ϖ�����be������I	W,�e�He���o�N\|Æ�����*C����U8kz���ǿ|��~�o��w�I~hh��^
	��N�*C��<p��)P�20l�aR7�6���'���*-�*����DWɡ~s��:\JFIW��g��T�%���Lq|)�lk��ce��X��C��}����0~�d�-&��N��S�p�'�`H�U�gM(�������ɽO���2��z��@h�`\�?�M!�c��1$V$'��e`'���4�_)�m�������	���=�V������>��ϯ]����u�P#�Β�P���.q=I>+��b��L*�*$
�Q���HLEfԊ3�y���L�X�6�k����s���q)���o��F���3?�*Ӎ����s�_��kǮ���Ύ��q�ښ�渃�w�h�G>S�:TC&��R�vIͤP�0�
�j��4�X�Og� J~|2N-�^l�m@g[뎭[ּ�v�~�LF���M)��"9.�5�rc���_�2|��R4���7��b�{ݺu��pMx����<-wK�K�qȶ�5�b9>>��y�R,F�E*P�C��d:Qq����~�g�����і���;gQQ����[vX�z�R2�zE��&�N�3��B&��.7�<�@c�5��\�щ}k
�k�)ګ�K4�E��JM�@5ێLn�$��$�I}u�Q������˹����`�J����[�U��5"t�dm��je�IyEk�����<S<��V�x��>��K��QP��<̌�<���%�t6�X%ѐ;$�(�F���={�>�LS�b�uJ��/i��q��:���P$�d$S9�7�b��}���I

��Z���a�	H[����+t/]�4
�4�l߹=�"����	��D"Q����L�i�R��x}n�wE��K(��zAmh��91o8��[~�Z�఺��$d8�R�q����ljj��#��#�Ǹ5٫9M'`?�k����Gǡ��"�^�z4���F�cTC�&28Nel�䂒9��.�����J�X��TSU Ĝ],�����˽^J�:E���'F�+�Q��S��"�������ō(�!�@�B�/Ћ=3f�"��'�5�Z�!�.��g
����3gΤ�gm-nv��2887R}����9s�a��$��Bt	�h5�(�U�
����/P�tA9���]�6p󢀠Y�A�8�b��<��"U���7ף:\'��IhEt��%~�8u%�7�R�OF8%7+�?��z�%��Z�'��E#T_�^Jjz]�W�TpԘ�V��)',��K�'n�>J���o��k��"o�������|񆺆\HA�!�j^�I�M�Q�cb��0H,`|b0�'�M+�=��S���҉	%��0sj"����B���	
������b�O�dF� B�32XW)5���NU�]9��+'��z	k���=�N�:9��Epr0����s�Ν+!	�b��ϕ�[�z�&�t����t�!L^4���P1A&P](t�x��&�Fe��R%.�ff�S���^N�쟇�.HW@��&��dw�ĩ`w�2�:�@�G��I��,�.._-�&a�Y�i�S�����"Hg`�����*�8A��ؤiS::��N�g3%Gon�"QlXsS�AM8��T22�4D����cg?��*�c�@��x��������pM��.Oj4�xI#<K��(R��'O�T�P!.�U�R�-��"H���A��T����.A5,�գ�ylx��r�R>���|��X&�"�ͭ"��� sl�VZ�N6�V˕�
�z<�R�T�'�Gvٟ�E��88ʞ��ɨ��])@q@��h`��{�Y����S�z��SC�JY��[N�8����?�S-�]������0�')ME�u�cPA��0�H���G�����"�t���ښ�9�f��aMw����懖�{�Ru���J�Ǹ�<�]F���aD�I|�OT2��ѐ�-Y+�J�i`&�C�p֒��L^W:e. ���d���C~O+����P8'Ii �������*m6�-���Xv���f��Ƥ��QX@�0�Ld$�K�4.U|x��(�I����J�?�r��-u3�A=�lx$�i5uu�w�hjm���Q��E��B~�Ո
��=��MMp*2�<�x���Ty��ƃ��Υ�	�oϾ=z��Q]pF&8�� ��b[��K��v):����s*S��FVc�guc�)}&��#�+��\�������#���zAy9�T:t�~�D��W��硳�V*��:qT�N���[�%nI�eF�(�p�:�x��4��1M%qI�^>Es�2S��D�E%&,�A���aL�el�X�r/��C?��H��E6���ƍ�L�roooSs�� 5^�Wɡք_���S�Z�/_�i�&aߑyB�*�d��݀����+�/d�h��֭[��-[�(L4��Ev�u�S����?~�h�$��VE��-AZ"vP�$�C��b�-T�!�4����ko�"(��*��	�6 Э~���w���Ҩx�>���ig>�d�� ��1��SM>�呯�!]j�=�~�� �"}op�3�FJ�����@ҸE�/>�Մ��V	.td��H�넦��!���������LL�s�.$�b{�|헓���%.7T{��c---7톏>�h������{�d����:o� �JM$�y`w׼����r2�mR��JEϮBj�ç4b׽W�.@�bi\����0�`k�<�Ŭ�V�0l������r��*,� d�9�Q�o 0/�R��#R-�U<4s�[m,[<B�
���t���fӜ�0�
���+'M@\�es��*,�ϴ�S�������H:�L$�o\�5�<����>B�`Wg��+S�0�vipx�e�����"�M`�3	s��U�����y�Qn�D�P�������nim��X���+.�b��|���ֶ������3�Iѱ�d0��锨taa�a�pg�y��8S>�p��=Sz�~�������o��!��D��t�s��"�)�Q[,6��5�cɻ���uH );�_��|�B��ߙ�v�pNԩ�	*�v0�bv�L
�4uh������;*M&բ������-�З�P�Y>�U����`�/sp�#���CQ�\Q�+*�*<YZ�Y�X\P��}����%�د����I�=<��c�~睻�;<�����?GM�\�������W���_yѹ�K]t�7��ή]���k����.L�xW[\/���Nȧb����9��	(��M��
�	���t{�.��0��x����s�l*�5�C�ӊ�2�5�����q� C�F!e�����6�a�MX"�U���|�j�d�*9�\F�)j�p8B�ހ_&�p�ߑ&z��t*+10q �bXͥhhD�楱��6~	�є4&�p+&4)1ʌOP�:-Vxk�xئY�
�>�N�"G0*�[7�p �aO��I�`�/���O=v뭷�D\��?��+X���Wtg�f��
���_X�G}������7\�5I�Sq�[��J��A��+���)�����'�NO�i�y�NŃ��1��Fs+)�ΐ!-�I�p�|��`���Xd�狜�-R�G:OĴ�ZI+�ͽj%�h������ȩJsd�* ��*��=�=Yҫ�k&S]��^3¡�y���<>)YBO�[�s)l+�EJ���@7��+�����.��jC!�p7�7��w�y�uZ�pJ1���b)�W�9v���v�C#�����{�654�P�� ~���-���D�v!g(�ϴ�5a�M�.�bѰ��2ɱ|!����<\ln�d2������}7�r��E+�<?̦��4`���r����Da?��xxp��H�Dj���!X챱@)B�D�'��]Ptj<�YE2��q�MsX̰&�CCE��%��U�f(T"� *�w�&y;>_ ߎ�;y���޻y��h4|��gO�bP:���s�vv�)�x�b8��Bϔ�TL&�KK �S����6n�-��-*�nJ"�t�q;��ʤi/M8"\G�����r��1������������%�w�X<�D,����Ҁ?�J����/@'6��y��/~�[jPu|\����8�B*���"�aO�Ncc�N]�Y&�ґJ5���\�_l�k�ص4�)�.O�:`
�,@���)�z��Q�z��[��-�B^�jX7���Άh��c�E��Z儬t7W�BL���+�o]��#���u�L6ǖDv�iRCb?�>�~mN@������gy�F���c���U�_{��84o��楗^j���"Y �x��[������\�[v��I����o��^�+V|���<9��K�MbI��r�<RB)*�]���\ N瞿T��w�1kꜱq���� /|����ɧ���)Ya|c4L� �/Mղ����ۯ�D�����R����F��K�]�ˉ'Fg]x(*M���&IPYi��r��B�J����� ͞=����ԩ��1��\&sŕW~�/�8��'S��B��ʕ+�@��\����;::�T������2s^��2jU�`U��J�]\\�[O���n@���]�P���A
�'�P}��8�V����XaE�Nub6�m�;w��2�����c�� wi�3Tq�yW��x�$�W{;9��TI��2LwK~V��C�|\dC�!�8 �x�GO<�f�x�d�E��!��D6.rDe�~�X�U�E��E�����b"1A43�_w�hA�	<v���=:N4��=�I*�����4 �x����4J-����GG��ZG��+A|ι�G:r��������(drCC�7,���m��<�'�7�Ea� �e�g������`�>w�g�zG���|��hM8��ǡ��̐ϫ;Eb�t�J�@eCٔ�	i�*��K��<�ήv����)���x�����&s�t���w���ӧO�`���B ��$"5�| �|㣀� ����=3  ��^�{���0)�[��`j3I��T�C�Nt��/F�T�I��:[�K E6�E9$M�(7k����Q���� ��w�lhl�j�#���Asi���ب���S�̌�pԄX�P���$'���Ԟ��6$� B���9��u�@�Ղ��f~�ᇬ�)k�PmH����������%�0�'��u{lr@D�]T�u�^=��w�'��!O#������C5��O1��j�c����o�4r����2c�f>%�P�ˮ�Dq4���^�p�;FG�[ZZ C�.��ttt��
����H�z0�cj;&�]�����	���#7[T�0|`|�V'���0v�����mx߾�=�%��SD��L�>�����Q�����8���YvThBc!hд�7x �$%^ʽ�ă�YRa��_=g�����_���ֆW���a��A�~NRI���=�ܫ��z߿��λ���m�}�'�d:G���^|����yz��|֊��Ɣ� )x���vh��g`y�l�x	��2�S���^1X�C��/�=s��ߎ�����S�[.
�N�GXzm9�tK6ei�*��Qz�[.��L|Ez��i�9ϋMe)s"o+��}!"���6TO�����-8a0��t+/Ԓu�L�օ��L\�I&�!�.�!%QaT��:	0��--����+�O�7w��ug���w߅݃Ҥ����	�
r#�Uу��*�KS�4�a��~/�AJ2�$R�422^T�P.�9<<���W=m)N$&��i<9K������2�,H��aLە mk��ᖶ��V)H�:���������<>�zx�,hh����|�tA�y�c�Ӟ�7w6�>	?����z����~������?w�L���PqU8B�}����k��𪫮okh����U�V���?�T��}�)܅m2�<v��;�MA������j5�9ԉCS�}.�ytp��G�G���C/�]+N>}M��,��w6�?x�?��^����g^x��> ���D(h*���Y�p��"L�)9U���A�PJ�BJ�����J2?�{�\�&VXGϦipj.��	�`*�ᾉ�s�W5%S�˷�YKޔ7�S�,!.0������h�/�$T��S��-��_���P
G��C��rK��S&!���Tlؑt�GEس;  ��IDAT��Ӛ��u��qPz�K�A���a�"���EM��i���O���]%M��8.�X�	d�W�����F'�ڠ
Ir�x���DR8�p��~c�K.zV4��*3���3�g�5�fu�]��w��@7X̘.���I��ǀ�������-��A(���A�gr�J��,,��[P�-��E�h)���E����\Z�>�����yc�U�#0qI �h&bc0�8`8��grr�N&u��6��b�P�7�Ds�mb�s���٤��}g=�9���ǳc�?v�hZ�
��J����2��Lv�0ŒjYx���l�<� @\԰�k�����r�DD!�x�e�/���v����g?�ӓOM�6�������.�		�W^���N? ��2o�<�k�����M�����̭b���`Y	�O���� Wn`�`�=��^�U������b1@<\�xuݺuC-��@���v�w8묳BA�|�M�p���|�}����|?T��=����qd�f!�8i'p?���f�1\^bS}���L���R�\��:t�y
ْ3����u���w�u�]����;qR�\�P��o�u-2�Vc>o�seT����+r���D�#������c'����#����-��whv1�kT�Ƶud+� �ى�#��TF�y�GqFDc�ζNYahfyP����Y�d�қ_dz�)��瘘�dR�|^�ILNV�=}��#CT�9�J�?SQ�gadl¹�h���V�%��x"f3s�-I|���"hB������U	�Т�>@&���f�)I)aǷg�DB�`��K�N����5h/�{{{wl]�m۶����UV�T?<�����s��7:6y��/^���-ZX�6OKlkk9yb0OÙy�'Z�Za�4#����<��P�b�0k4��w���҅����{�@�i�Ʋe�>x�jA�q`����LUd$�J�<��E��GI��:��Q ��BX:p�BJ�
5~/v���7�E6E���dO��P(�t��\6�x�xdl�h����h�0|arY�����S�d�[�m��2�;e�E �����]��BMr�*6���m�����~_�&���R�l]]= ���	�L���CUӼ����d["�Z
��Nsҩz��9I���$���D���/���M%O���=�O�(
ꥶ�8g��A�%�yp�X(�O&�MDK$�ة�*TJ�J�P�#M�2$N���B^T��R[w��������m��OL�m���u�P0���cC����Ի�8��9͡�gc#��<�N���<jgg���i��>�$��7c���sE�d�jj�k"�\�@іŃ�\�\4+E�y�D������r6��Z3Ceq-'��c=�Ӱ�.�'�Κ�2��4���}@>�5E�+�.;���ϟI'�p����:gΜ�S:g�^�ࣂ���"�B3����h�S8w�����w��a�S��R�x��x<òp��i=�x�\詧��[�i.\"G%�
۷T:
�n�����dM4Rb=<u�����d�/��;�2�G���i)W����Ŕ�x��%p\��"4~=��Y�?̓_�m��҉/!D�A{�
�{__߁`�Tf�.���M֛�qrRԇfz���ȁ���sm����By;A����n%!w�|%�d������d�>U�~`�/�#ZY�����D�	���0Dp����(פ�+q�/59�,�Ӵ����̘1#��g灆&'�mZ��+�t�<���Ţ]�s�A��*E
9�����ƃ%��ͫ��}/���@ᝆ��
!�E�Đ�9��a�<HK"K$O$T�\���7K�[L�9�J��Ì5���]!M�ݔȼLQƳx�ּ{j'������,��]���˗Cd�y��b[�Z�MܣQ������/����ol�uD柒���� �?�{���҅�o߾?�g߾=���?��˯��A���34��{����:ٹ@�t7\;ݰo��5/�
Q�1UR��ǎ�r�h�����vj�߉ !�ΩF��U���o��3Q��=�hmm�c��~ನߕ�d�(�3O`Eۛj{O�A��g�S��
Pj�p �F6�[��魵@�c	
]X.���T�"n�`�S�U˃VH/�rv8λ��+:>�d'b9+�����X����X��t�|���sՊ K��=[��t:.�d~"	�L���㏤Λ����]�*G:���uXb�|X�u�Xl��1�\>���h�\����UC2:�"�vP���/�Nނw尶*�`����|�b��V�����(������Q����.Z�����8�!��n�;�p�&Kd94��|�B��p��١�̆��tM{}�FE�ts�"����K��8	䕹6b����L���gGiQ�4I�����I��eV2t��Q*�����([`�(0�������\A�'vy=č"HgOfE��n�X�Q�+����K/����;w���������/�ҝ>�`��ڠ��0W�Y0�S�,���;u��?�7 G�J�u&�ƻ?��<r�ps<�bŊ%K���[�*P�	{u5�>���o��O~��4a�%Ϧ�4��]����\�u������Z�͙��3g:܂���̓)��"����V�0���WO;�4n�_���{<8��=�81��4��t�޲eK�����NN$�M�.U�}�^�7eʔ�����Ə0��s|Ήޣ�]~9�`m�u�K�%����FsyB�N)i)���Z�Q�b���U,*%�Q9��y�7͓��0s��Y��L��Ei���5�a�HH]:t�9Ѹ׮�^n�""�-5_�V��GΨ��GF&���*�����aVse�gJu��n
,�$�ʍ
�y��]��J�` ��������9	�J��V�
,�'�F��0��AjЫ��4�D!�,FXl�].ZW��C�qcu�-̉V�\�3:��.H����\1�[��p�JLD$�!��~��?��>�����Tu���ׁ8�mK�,��~|�w�;S�N��A��k�⑏�U�d���nx�;�����~N1(e�N�;\FkG�D|7�b�X�wG[�c�����UgZ�h��kɒPH*��D�V�#j�uS�@p]]],5	Q9t�zY�C�^���k��)����zuT.��z*n�oh����~헎.Z� 
�|���5�x^7N���.���K����O����V&GƟ|�I����~8�~C��HQ��������X19>:�6����+>�^.Oe+}}'�7E��x�D���ި����Ϗբ�L�e���b�"��W���T����G���ȤN�m|�㠛��{������+)����֐�'yI�ׅ�%���2�1U�%Ё3���0�uJB�o���;���WiSz��.���v(S��\mJw�����]���A�-ȳ��"e�Ir����-~	$U�'w�>sR�А���ں��V���(W@�H96��j9�(������W*F(�O�Y�b�$� J���S��er�;G!	HV�*Y�ʃs����ՙ9
��)��4��[�Y�D���D�n��y�F���t�-B�B|�mm���|!��h霿��/��ac-aϜ9+��C�iMuF�F����_xA"��/[���3v�D�szfJgkWWp*�P�R�v:-zE�ٱ�555�Z�|� �L�U�ǣG�P-�����E���Z�����g�����:K�#�Qi޾e����0��O�*����*ҫ.����g+�7�+>������ �UOO7�z7�Q�Խi|,����� �@�P��!ط�	[)ӳ��[:��^��S���m۶Q��'v�矕�m	���H}�HM1����6/.������"�;/�Ax}��ex��$]��9�������|�'�wpuQ�����MB�˓��"�=�ϗ�|�$�TQ�\Qe���x'U�pZ���%c� E��a��(��֘�[+le�.�F|y\k�g������ a�h�&w���J��Ra�� ^Go�w�o��� T�T����z�S�R�hF5� �?a���|zjG�&2ɣ�t�~������s�����8�P}M ��i����z��Voltׇ,@ {���w,v��+����q��Ǩ�['�$��`��Qh���Pè�����Ǟɥ�^��Ά��n&���!~6�6�����ⷉ&Oٻw��W_��߸��_�`�8a� `!��;�܃�}�'��V�Z�{�[������I�.	Sgj��ipun9���Ո����؎��&��	�K������^���-Y�h��D(�O$c�-M��B�eI���9e����8���Sajk�ݾ������50x��կx=^8�#c#Ϭ��������pdl���j�
�h(/��pķc��L��H�!?����a�j�u<ǻ��������&Dݾsǻￏ32��=��O�)�(9��vI%6׼ԸKBBl~�q�RIJ\�
��-Б���K[�`?��$�'�8�/���n�7�Ũ�i2IM^A���T/�����	d�T�Z�"Ǡ��d]�؟H�T�lQ}M��V"Z~��E�%�ƪ�P��ϯrY��$�4`��
U��9
T�͜�L��J"AJ��uB��N�)�19���ʎbK���0��D'J��c�:5��?��ȑ#�g����w�_��Ï�ٰa������b>��!�2!�b	���%����5wwuus�Q��mh�o�Y�wQ�o�Ɓ�2N�2D-Δ�x�h$�����g�qF*� 
ۅs����׵�!+d��_;�b��l"�[��"p0�������y!x���o�m"{6�/�� �qy��^�iҝ��Aá�M���͸a����Ӧ��H���d���Q�&C�c<)�k��1c�����"4@� ���݋�N�~�k���w+%��N%����bG8W(@�#{J��IV��(���'O�$��""Cf��L�>o��p�=.7�7^��twcM<�>	_�`]����V�+G)D�,7��]NWV�b:�zt\A�5��Cn�V�"IA.��+�Vܡ�0�@�,����]y��$!+x8�o3ϊL ���5�2�FJ�+DN���4��ή�0*���J��JA�*�����+?��8��J�V&7V���������!R��g�]}��W��Q��G���߾�ꫯ�江�R��b�Őda�pZ ql�^|��~�{�⅓cc�O>���6���Y�	��K�dE#!.�+GG�=TŨ[7o��7�7AGZy���-(˛N��n�O��L�gŜ{����F~�4�宸�W^y�_���ի�{466���WK�\.��������Μ�{��pMnU*�inj�T���#�/�M����fMs�U���4�����1�`}���*.�769z��}h�A���S�mٳ�øuQ�^i�ĎQ�a>S�;{�t�W�G�Ǆۦ�8XEMq
LN��j0�L�YP���ӧ́o��l|�sc8��-��*'��ݺk�> N��pwO�Ёg}g�{�O�S;�:�����e)m������M�%؉��2�d���.���u��eQT�`����Ő��3>�~�W��P@��u��,�:y��z�FE��L��I/�
��c���99��t�hQ���o�@�jB�\ⅺ�vH�l�T�T�����hՐ�/���(iy'3�˸L���%�[P��{Rb�Z)�Е
�S���H���	ܷI�)�-`��Q�GU`i8&�y�_�]�v�v�W׮]�C���\��O��W^W&��Rvtv��R����!��Z�I|���e��G�c�Ǉ�!,�|���@C2���M��J�2Ễ\<�zϞ=8�p�֭[��{q+͍$�4G%s�(�����D�$$֓O>Y_e@&4�T���dՅ�~��������_�����ӊ+p��=$i�j�L�.�Hy�2��3��̉�����}��_��յkayBa}d��:eQ\�k�ҭ[��75,[���CT^T[pH%�^M��_�~ڂy�ãu!���%�9�۟H�{.>����JT2��$�A|�T<Au� ���g@�����nv�ut��d�-[6�8q���__�hQ��:��%�{�7L�*v��)R�'i<�P���X
Vg�P�ф�k钺܂Nﴝ�V�3)�B~���%NXf����J|��	%�)c@=<�m<F��⺔(+�.rdR��rc�u�}��A1{��Z\���"��tqn�sdH�����je��X���(�K�,�Va��ԲId�\��L+��}ª�}ҜV�h�$��<��"�N�=(�Dt�_�yf�����w��omm��$�Y�-),q�� (��a�傁��̛7�k��|�M A�Ϧڠ�.2�`�v׶-R�.9F�h|lz���_�������� l�]��}����L��^��+����h骱f͚m�v�Z�4�v��)OM"&�F��<�ѽ�>���n�|o��T)�?>�����Fd:�i��|��:�my���||��B��ǒG����#8=S�ñܵw>;�{J��c�LF��㭇ּ��gK�z�rY���|j2�?:1�K%�ť�ۈ��"���:����2n�\�ԅ'���&�yKk+��.[��KV������ܺg��+k_ݿ� |��,���94��j��޽`����v��+�h=tЋ{ۖHN�������3�PH�͑�q&�wC�Id.C�5��C�(��z~�CR $T4^�e��^&�ue�9M�`���a6*_@0	OR��I$��A[���L�T��SS��
�C#�UG��3����:iwGZEB*��R��������`�ML&u�g˃�9��s(�����A63�<�Ю�Lt�bgi��P�TJ+�#�c��nHD�ld�iR��H�(v���r[]���������'S�=�"O�k
Q�>|��os��7������4�3ѩG^*J�N}'v��:�������M�-������K�]s�yX���Ý����9%��h�ε�+qOd7
�#Z�r莭[������ŋ��b�|󍷾��o�cA*q+�^��LϏ��������/^}�%�pS��>v��i�I��R&5,��K��w|�g:��x �+W.�淾��_�Br�[i������¦�k�X�Њ'�\�Z�BA!��d&ZW7��bS�B���{�w�{�
��4�+C�y��J
ݹ8NH���Syq���^JT:���ٳ��?�a:��*�x�%���dm���s��-Z6�����M�,Wt�i%�_bK	Sb�����OyN*z�hH���6jb��-����U�����v��d2�{vSk��<¶�TfLqk��Ӡ�xI�Z�4�(�4<��x�{�ާ�DNEȀ[��lR�r�$��ID�T��7��W�c<Rc��U�$��W�ϗ�u����E��Y]�J
ل� �S���O���X�&U�҇�����%J��`v�;�Q�gׯ_�q�ƳO?+��ފ�	E	_��IB��b�1MO�Z�j�⥷�~{1���{�h(Z���p������K/�D19MH�iR/Q��ܮx.��^��u�lP��K.>}��+�.���E�%ꌬ�Bze�+�_����YJ�cY*��=���{xU�p��C_���>��O�&�>����M2[�	2LC/�Z����grT��3�{px����'�hmmŉ�ꪫ�}��o�����ęSؤTh��P����,��a�`0LU�)�c�]z�3g�\u�55.�D��޸n�aFR��"�R6	t��if$�$U��tӍmS}�l
�Ǌ�+��E	hQ3�'WP���&�26�ܸ�#�< �%}g�<�<��q��(M�L$��)R�Rm�ӥ�c�����q�և7���<|�|b���jpx�pTx֬@8�oߞ|&C���FY`,N�4���~�acE<\��3{Nl|Ls�''�$����r�>'Xֆ`�B����f��ti�c�D�lV���9ӕd��	.26:Fw^�A���	�^qd�e�)����9�2��?cBRȮi��1�P0Hڟ�?)[�F�߯��#�gU���e�������qO��ڏ�dΜYX��>���p��ln��]�u/������L��	8�8�����3�V&�Z�JvNQo�wO���U�;hz��b
��D���T}�\u��ms���}�ɦoz�B�A���QA|b����A��SDP���A�H'���4ҳ��f����>wn��93#o?|���̝_9�|�k�ᡧ�~�f͚#�-�܍�cӧOw��/�������kJ7��>a��3;,�N?��#}����P���g�QC�����6*1nqx�ze�$��QM�6<g�<�������_��'�q���y�p�$��Q�.��K4�CL*��szݧi����b��?����7]{��Ep}��^#K*�X��Ysq�Sy
�O��g�=�����CC���9�`AW4FLR�.�>F�8F�B����2�V�0��Ys��b)jZ��`gE��+�)EHX��- e:�htr���R�\�
�Ĝ�ˋ�+�+c�i���%	?b���cÇ���Vph,�qs`�>!C{y:vǙ�$�]}�?�h���ԙ�In�R����ƚ6$�mj�)�]��$hj���I©���Bt��c�_��������VQ�H&�� �E��(�{<�G��Zaj}b��k����̨�a�4��j���14Q��]�4�b��%o%�0�R�7I�u�:餓fuw��Z�S��{U��Ν;�x��^z���z,8@��b+�꡾�H&�)���������ٺ3��H<f1�����[����nʔ`����\�Jf�*�E��|���^��S A,>�H����������90�����19�=�c���8M��0�]��F��/��ں�����V����o�}��g�u�Đd��0���`#c�r�J2-B7hH[4
N���ĕ<�ԓ�mP��v�x埯���?\��eҠ],����B9�P��ϩ���?!��w�O�:=m��=ok������AJ�s�x�@����a�U*��[tyO<�&
x��U��BC@|���
I���גP2�����q�YgAJ�(��ޞ��T�L2��˸�x,Zuj]� П\�38�ӳLJ��3Tu�5j;�{ծ��p V��<|���T73��Z���4��e�nZٜ�ś�g8�P�<党c�dȣ,Q�|���I�J�C�U�����渱T���|��ј1<2eh	j#P�R��k��Q��a��Sv�ʁ��m�x�.T��U���q�P���\!O��w�s�f���&���R�
���TK>�VT���K�Bz�b;VHX�`�tF������.�(x3�6�͔b��J��������]n����?��T~k�w_��ݳ{f����	jt�(��]���}87V�;�Q,�kNJ's�39^}p� =�w!R
���7��i�:��6�	�x;�=��fTj�.� �9���),1>5.���쒔�jSG�z����e^b��7��g	f	�+����N%�y�����x�"Eب��';�Z��䃝�R�>mz\���փ��7���?锓qg�-�povm�N �ԥBӎ���M�q�v�m��fJ�b7�|�G) a�G�Q��l��4]�:�݃���9GxY�_$Q�)� bȡ2����A�$̃yq�pp��vQ��I�0�(^�r�J����{� 	ҡ�!ԦM��XjO>lE�+��� �S��]��C@x6Ul�aR�n�$Қ'@X��/<�Vfo��"׋��v�.4�	RVAUҺIQ�b���;Z�KR��M�H���9A�ÎY�@�rJ̓2��!PF�q� ٍ�#c9���g|;e�P�ZZ�9<�A]]m̽	�Z�O��_�Ez�:�O�L�,SL�?�J��H���u:�W��0�VP`�t�'�9E���F}��IRea��f,N�d���̖�i�!<��)��)�8v.A�
��fHB�`�OFZ2iZVK[kٮ��-m#b j���I����Ѩ	��#�I7s��+��]��+I0���P�Q+� �㉽O�)hF����Ɉ�ÉMKv�4ur�w�y��uT'�z4XFW���X��O�>}ޢexN��5�;�wC����_�R�:k���G�X��Z%��6�{x�!Q��;�A�%&t��ٳ#�m�v,\�vH̕KP���~���ҹՒg�@\A���o�ꈧ�Zu�D	ȋ]�=�u~��Kv���i�T�]bn߾=ٜ�ߦqNTLO�b��uML�Dss�.({��-�	�C1��	i�<�*j�C�3�ʅ����p��C*Tx�2�A"`�����.tr��9�!�\C�$��ZՓJ#(��c��S2��aʤ0��7f��#�TT���/�L(�'q�F|��H�(�Y) ����ݤܫ�E�q�l����"\q��P$Jc��!Κ2�p`
����@]Ij����Z�FW��P�(n��qW�$���ɒ!5��H0	� ���e/@��Cr�D{�����ጠ�6AQ5�āu�-'y��L��4:J�$U%�DS~*+ڃ�gP�ǰ�%j ��Nu0�$��W<�J�Q�X�NL�ܹSa'J�{QF�QX�BE02'�a�+n5��d�pt�A�`�4�&/�|��\(B�&��xJ���-EoU��H����m�J�Z[d���s:���-�7�<��*�ZZ� ��P�	xx�{aJ���:d��=����w�b ��*����3(�/.d�Paq��Ӧ�m��"X��g�yf,���r�"t�D�`� L��ƭΙ3G�={��`�?w:�5�;�ꫯƣ�4�5\k� :�|�d/$x���e�Yͪ�h蚌��,�$hV�OUX��P$���l<YL��$T>49���d�1!yWJn��hQeˍf*��	�W��C�P�#n�;4���p+VF�����@�h�{���|����Tˠ� _�7;��RΘ�{�L:��C��84\u�"��˧~pҊ����2t�=(5DBҵI%������p��3��"U[��Z��ǅ�1�v������rB�u��"�r��5�lLӪ��,$d����r.��MNd���_a�m߾�q�'>���GÔ�xo᲏@�l޶}N��9��	Sӵ���!�0�[[�A��Ǔ�ze�,)A�;��!vո '�{!rT�Z�͘� 6}|�#��h���V�)���L�N��)������͙������N�d*~��F�e��	��d��Uv�|z���W�d%�4�D:��iQp�uI?��ċ���V�t�=�t�*�k�Z�Ja�	� ��^�@�������-9����SWљ�H�[���<�)1I�_�r8J��p�����#")AE�6�BAl*��*�)-���9��ö��R�W���<&�Z���ZYi��KX�qq����;O���<5����	���܊����p�P��0yؙ1��&�����ށ��vClk1~�������:<�$����]���xL��zv�Y��L;�h^������2�Kd��UQ��� !7�d�pA�%[��}}Iga��3�!���KaBao���4�} �*;`��M�J<����@nl�λ���>O�hhr��L�6Ңl�L���I��� Q��}��C�Q�+�|��K/�4�&�[�e7J�ay�|H�J��m�_���mH�x�!��5%BzL�
V�q&���K��3f�w-� 2��S"�:�ʺ
ki5��{�D�1��˥Y���j���o���e6���;��5�"1O]�
(�3�������l�0``�񏿓�W5��^��q)�Z��Z#'!�5t��h6ڻ�U��]��B ���V��`��l�bU�_u��{5l�Qt�1�R��G1(&�r}N�)]�ILO�d��v�.���tK��0�R�M�靝�a�
kV�W3 �b�����T*�b�2�V	���H|5İ�)/V��*%��+�[2�eW%�������N��FϨ��x&�~l@�rE�*�N�X�$a)��������l`|���'���y����*��ƴ��NشjR�Ό����p'��/\z�y睷���{D��E����k*Jx>N@�f�#%Ç�Ν[���Xђ%K���}���ڽ��[/��$;}�܁K�\�҈��*!�ҢR �r�[��]1��/%��σ�L��Z�e�̙'���0CTEy�̡C�@*4�)��&�6�%>�R���%����c2�rs�en)~))86�T���(�ڱ�M\��g�����{w�~��W����*��u�^����A�|D����c�T�z�MmP�{v�򱓏���b��ܤX!���[�;ĤOKЎZ��^���Aab{#��'�f��O��H�w�F|Őj�:ˑ�s��m\5��Y�_�4|Q�C_f�Q)�
Gb�.j���K�t2�9�*�On��@`�P�xX1x�h�^Ȅy PM��*W�QO�q�)�����=�*BD�� iit#�Dbȫ����6�Ӷ�]��u�P��p����kE�,�V�k�D���<�&�$��Qf 1v0͙)U�A�
����bZr�ƮTd�3��<W�*� l����k�������I
�,>�@4��R�;	��;q�A=���7o��(E}�p˭�\s��m��y�t&#ꈤ#� ��D�%T�%�bU�7���7�+K|q��x�t��˲\"QP)�Y�_P�y̰�9�s�6
J��{q��ʍf����V�f�����Vbu!��A��5�^�T���9���
/yUᰂ��m���39N��-x=�>�،��+
@�(�-3q��%R�x���Q	�5���eC_��2�3j%�Ҹeq1j�>����G�%Tٲ�H�d}�R
>��!;3�R޲_%ªh�_�U߯���Ǘ_T��y�]�Q���$�������pJs�������qC�P��gW�t$�Λフ�%"S=Q��b	������P�^(�hF��n$b���1��xoo����9�|��뮓�U��ݸ�nx��W�RTW����i�ny��*s�C���ha�C{��(��0D�*�j��:)�f��d\�0@���i /��6��$�WzO(32rꩧ���y��Șjj-���}z>���R!٬�J6���Y3f^y|ܦ��U�����wu��۳g�[.��E���{n�XND�^'(
�8j����^J�R��ij��j���
Y�jՖ-[�������L(�::S��$7�;��y�8pO1�,_֚̕bIw���+Va��z�8�7���{�M�ϟ���w�'~���~��_����)��j�ީ�p��$��-�����N���k8݋.��?�A_/���r�j<�/z�4ӂ��q���{!̟�yӦs?�Ex�C�H*_?��*�W}n%oL����{�\���6.,+�?�إҹ���oS��ё�͌��.�\dfؒ��,�Id2қ&�&��Z��n��4�8d�6����'��))#h����WJ,������?�iû��̙�F�ra�2T�z����X�;�*U�p�pH����M���"\��8f&���LC�
�(@o��B�\������R����W�x�1�<~��?��� SE�I�OĹ��1�R�S���L�S|hN"�׆a%�����=:z6���@3�e�!����Un����	�iTYc��Ϝ�O}ꏷ��9��O�D�:�d3I��KLrꙟ���~w���;３d/ƮҲ-�E�v�F0�W}��@#v��2��|�J�U�"$�q����m���ׯ���Zs��3N;�.Z�n��#�:餓�;��_��W;w�����}�=�������`h�o��&p�W����Tr��姝v��ç{�r��g���߶m��U0.����m�reo8J��`�*�H���x�P3`��z����!�v�������D�����Ϟ{�TR��>jYRВ�Ò��Z��K�-$�*�N��Qk��ɲ�	�a��R+��������x�F���ǆ�)L��kq�֬�(�I7U��[��� !�Ԫ��vs�-=3����%d�E��Rزy���LN�|H��"-����&{�򐖞��A�}�z�|�(�I%����%3�D���f�ѵ���	�ߵ}ǚ5k��^�W���W^y%�Jb�W^y�Y���}�ݗ_z�g�	^��!�Fd��0 څu���>ƹ5�#cc��E�C��@�5T!����ubn`X����=sf[K+�vU�A��Y<>fE��DaZ�ݽ�Z,}��O8�+�q9����~r`��?8������oh`���Ϝs�̙3��.��� ��^^kfdb��6�=�FH�L�%
4ID��y�I�@ݹ6�K�(����y��۶wL�vх��ٹm�։�	h���?��^�P&�o���[#�d�O~��j8��o���.�����DbŊ`Nl�}������.ϴ�������޾���~��K����O~����]�x/|N�2���x,��E(ᐦ�k��_�s�p��������Ν��&�����-�����6��.�m���R����s����'�M�&q�$p%~#;�?��@�6TM:}v(�����s���W�r��ht=�n�Q�q�R�kP)�Bu�Q��D�؇%�H��q=�XkXa��!��V�%�I�.�Ӻ	ZڭTC={?f�����JB/��*�B˓�TKs��9��CĄ�I4dMu�}}�.8��3�X�/��k�� ��~��^�-Y���/�	�be�������x���[������ҋ���/B�7
���\
����s�tP���m�Fp�e��u�Y$)zzd�l�[b?��
2��`c���������s�='�����*6U��X���=�ؿ�v^&�(��P�+R�J��#4�/�2�ሱ$xϼ�*N	t����[�����TzE����`�[����aS�"jxJ}�����륩��e�ر���Â��ۼꪫ��vK3��������^~�e�G�\[�C$_����G]�n<^�A���W_}u��i�|�����~`� 	x�Tєl�N�rE� ��t.I�2�`;�d8~y�QG����4�G���7֮]{px
��*��H�3oΒ%K��T{Msi`��$��	�p56�b�taHIr�#Ĩ�����Q�6������|V�e�bF�w���(�Qf�7Ќ��	�Q��CA��_y2��/�6��$��q���,��RS&�����TWW��蘐PCo�b1Pj�=�oo�>��o~�
����)E0{--Mx�׾v�=��\s�O<qx�P,�%�AO`B�}�C�/q����i���?��-�܂C`򔓿��/\q��*Q��JU�`|����*�g�����~��4}�s�-]��g?��.X}�q��4p	VdR��*#s�t*�K���hع}tW��@���R�j��V���>�3����C�	r#Ǉ+�����-�d"U�9m����#�gs��)x���P�DXn9HaIظ	�#!(=��mx�M��$����G�.H�iK/ò��~�R��Z�`T�O<��?�
�	/�z�����<Q()�d��^}��p4���Λ�y��g�|�-�d[{��?�(���n����������Ǩ��g������)�q�����v�D���"B�x�X��X"���EŶ�mߞ<z弹=V8:9�����'� ���;����͢�o0+�����v�ϓ'5
@8�d��hOa��|�tE���xXE8R"r$���K�"E�T��S7h��V��.��y�Pʱ�F���YK��Tq`�2e"��(��gz.�6S	��]	�N� �@P� ~�Adk>z�g��ѕ����3������2��g��x�t�b���Nu*_(ہ���T�T>ys�'?�I!��ϐ�Ҥ	��#��D.������`�瞻�Z�
��4��	B:�+ANϚ=�K_�� �p�I`$/^�{�n�ب�Kn��7�R�ℂ.���"	{p)����;�lذ��]�T��W9������XIGk�׾����V	�R �\h�|����R�6m���|�=�+v2e��ip�p�8A������U�.U�����
�$��s��^��$_����H�7��H��e����G���,��T��=�(&�KQ���%���{���h�t/�(�O$�����O��ʅ�KwR&����3z�VCIҡa|2�������ө��	w4l�4=׷i������AB?�pS21>>	c��V�6�[�C|� =�qiT>eEɜIVP򙂔�"�#�x��Z������5[o�UY��An��j�� s���������j����,�f���{���|�y���
M�K�͘�	���_�,��?�x���u��Ac@Ön���2�^���}���}�������`�>�8�J�>��w����駞Z��hVk�)��K&����.)0��{�@��պ� l�t*Ei�: TpT��O��F��3��xƾ�@�0IsS��{� U��V�;�)�$e���b�/>�|[[�����|�,H�T��8b��54[+���߅�\��SR�ݻv�����F�eW�잣'��4}�u4j_l���o��S�s|xX�2�t�HQ�����i��2.'m�iUS�Q�4�-"!��+�[nin��s�n6�gZԪ����(M;�>bE��"v���t�r~�P���6��抅�e�`�I-��m�I�0pl*Mjj� :�a�I��r�Ga�
*,><��M�{d,_Ac�r��I8�����gy����].JE�'͚�#�:R4%bQ�˓Y��^���a�kiT`k�[$Xu)��|��H�F�ڇ���p��DvP~��UZ�K�(c�ja/���2�1Ģ�t����p,�<�S�~����Qi����ܾ���B|l��s��W^�X��T=��6�R�hN�8�c�.�я~t��0���w�}��I0&��aF���?0s�_���p����`p�tP���?�m��8���< ťq�Ňz�����X� �L+�*tk}���+�"$�V�")N�8p�:;!iʕ�	��4�XB�x �A]��6sfW���4v�+�:�Ta�
|�ƴ�$%�����ƛ�(!Y����oo�eN҈�u�����##-����6o��*�1H�V������Rǐ�D<B%N6�K*U���~0�J�e:9�>��$��Q5L�ۦ��R��'9I��E5ǜ�"GL/�H��@t]�7�kS��@��T��d�{����l�cjr��9i�d&�H�fa����05!�H5��P/��N��Q�n4���^���͐���84N�ɖ�x�m~��_�,`$dR�;e*���5R�L	"h5\SU����$�L!Sx�T8g�L���h��B5[&��b��8�;�8�� �{�
!�4x4N���y=���w@E[6�Պ�m��ҙ֐bz���-�Ԉ{x׎��ɱ�����#���.�0bq�Gq���Ͻ�+_�������H��.�/�}�W^��>�ۘ��;g�sϞ=7��ƍ7R���7�$&rvC`�֖����&��s����Ԯ��@�R��N�_D#��^���}�m;�V�jՍ��"���w����[ҳ�Vۻ��xvd����ԩt�dS�-p� ���	�jP�Djs����`O��i���}{��Ec$�FF �����r%���hQ=�*���p��Ri�mR�8�
Y� n�ï�c�\�Z y�O�_�}�7Y�29j�kj�?�54��V&�s4�&�r�Pv*OhqQ�m��
E�1lP��:�M{��!AR����t��M6��\
?Y�]5��?p`ќ�i�g���#�-�/�[:��K��}��t2U�	��BP�M��������������*--4"��S�}�9ѦhN*��t�0+�QۮF�i�u�uT�]*pj�}<
��J�u�pah�����L������|��S�"D7&Ѧr�P�)���APNB`ftE��J�G5ì0���a��Ԝ9�S�i� P�=�w��c��nn���*ە���/���%=s���_y����ەH��B�e¤;����8r�³V���[��͝6�p��8�bN�&��Pm�����ի�����{wc��#�`�D"�2�$yA@�/NM5��щo~�W_�pj�7C�J/�oWWW�9�_�M7��)&>Dd���ɩ���Td1��:.��b������]8p�U�A��NW^~��G~�d�֭x�xv\��B�8�A��K�b:]|<1{�?�J�5J��*a̸���mnJ��'�bS#�������\��j<��֤h��"\!��&�i2��\�P�D�$w�����x��U��tsS�����8�Y �p����dC7���VuE�^J�X5��a��.|ܰN�>��	>ꫯ��ȣG���?^y�
�0΅�R��b#�
k�x+<�8	K��uE�r4,
�R��س|{��i&�L�,v46b�,�51��W�;3W�z�r�Z",�E�U�+R M�'��#$�a�6�Ԛ�Zo�o���,���������G���}��8�X��=,M��ǯ��j�E[W;��F#N�p�	'��0p�5�A��)�=�a�^J璭�+�m�t�IO=�<N�#��Av�[���B��gA��2<�)��5s���ۆ��g͝�q���+V���i|S;�L(���T�P��X���5kΚ� ��]I����6�D�:�^աjz����UTa�Р����{���Ƣ�������Y��߻w�ʕ�����}8i+d�Nb1K3��%Un����ĵ��	x��#��ۄ_���ˍ�7�h�^�����b�I��`� ny���8��i�a��O�UC�*�4�R�2q�,U�f����D%!�e&��cq=>�	�����|���#q����!��y{������mCC���y!2O��\�ɭ�5����� \C�Q�M<��3vh,_����1XN�.�1��Ͱʸ�xx�R!>�)����.��a�]x.!��d��7gR4��j��NC�a��'z�c�U*�/��|ŵi܀�ل�P�h
%�Հ��}�H�  6�'E\�g<�D�&]��;����u�5w���`�Ǒ�(�'�|��)�˗�����AXs�f����>}���9��6�7{Μ���G�s�-��T��P����w/��<Jwy$��N����{f._���^?84��b%K�~�طt0p����e�8x	�  '8G�)��Z�<��u��� <�������{�L�3�~
�,)ٻw�_���ܺ��O2 �Wo�Q�HX�\���Z}�&��z�ZX����*ħS�#%�xWww7A��z}����|��0O*_���:�K/<��c���O����؟���y:����aZ|��������ɷtّ��>wp�����JC=[��D�Ze��%l�i۔���	�rߑ
!�2��
R^�]�3�#�{�wP��	�9���M��Ry�;kQ����qҤ�\�/�ԂH���\�TQ�f��g�8�=H�^�U�&n��n�'�K��w��WIk�4�ᄏ����7�5��o������l�2q���'���qnM	�!i%1�2-�4Q3�FrO��F}fC�7b�A�_X��S�5up	�rLi�kKWj�!Ŧ�Y%�NSS��W��cǶ�/�[8���������������/S��o��	Ʌ���8�-�x��i8
6��jn��e�78v9d�4��Q�zB���B!����KK�T�½�����}��r���o�G�dU��l�]-�L9�X� S��G>�ٳg���?�3{&����}��{�_�t+�h�V�b�� >��I|MȑYp�`D��{�����������L�4-�X����jVĨ�K�,�#AKd�	ʅg�:�<��R�����w�$	f�4���`]H�D,��3r۞y�o��cVAޛJe�qY�hngs����%K�,ZrdgG����X"U��#y.zR$���uF؂������0AB8�'e���&���x	^�� ����KCluB�h�?�l�"��0d&&Ƹ�ؒ��J�d��5�A�"�H5�WH4�X���
�lmN1��OU��::r�Kg憹x��72�`�I���O>�K_��Ҟe��xn,۰��W^yer2��_p������ ���:��~��'IVqZ�x*�:�T�O�E���a(gn+��2�Kj�C`ӈej�E#�\a!ips�`����*�]18��V�֩d (@U�=H`�ٷ66ON�	�ch`����|�+�Çp&��Y���O�
&��_���tB�&T��{v�랛�¥౳�i�|��?<2l�p4^,W[��؆ēJ��q�����c1}`�*�6mZ�2<:-P!�j�<%���ƥI�	�����ĩ��Ε����/�x㍯���Bm���{���v�FTN���_z}P�DҤ���g|��.Y���r7n���/7��&�hY�"��e��7�c�X��Bj-��C8��7���^г �ܾ�wւ!�Qʃ�F�,�N�m۶Q�{wbO*��y��yZeG�Ϛ3��O-bm;��.�d�������Y#Y�:�}�*i�����d��$�DG%�,'�!O��.
�[�X���16LM�����Bt&Eq��n��5�@?���/��q7�ʐ-T�>���!�mބ�Y���Ͼ�>h #L��6�� g���W����T��W��{�BP4�E���5E�t�ͤxEȃQ	MV�bB��a��kB�F����%���tx��ø�T���g?{�UW]u�%_���O�i Y%�{�ْ4�d���X̄U"������f�lMɌ��XP����́����{�=����r"I� ��[�c��UGO�箻�Т�������᱑�����NxXJ_�5�\s��/��>������χE
휝��~�i,�6��*0�A��A�j�\+�ѱhPo��$�[o�����86��С�w�}�����ǟ����k�ď8�o|����~�z4gZ�S<նa�� @ ��*��k�Y9(Qj��B8E��-[��2ݮcFc��N�v�j&�l�׶	�&>b��W_s۶f�^�y�9;u���Y=:�R��NL��ܧn��f����/�C���V}����`���8I��q�bͪ<<�����}�k����tϜ�DF����X���|�*Z�9��A0c�R�EM��M�R2��ȴ���W�^!d���[{�aO�aAQie���(i��{{z���8l�駟����<�.*B��5cLP�Rܵkk��{ �M-LC ܪ].V�<7��Lp�{l�[m( ����Ձ��͇
+�*�F�%%S�iX�n]qN�x���i0��r81MAf���I;�S�n�
^�Y@�e���veǎQ������ֻ�y:KQ�|�;�3pp �J�&)�p҉'r9�P���h�1�CL�����P��)����m�⚱ �>7�[c��GB���)�s6o޼sǎ�˖A�0� �2/�����+Ww�1.��A&�=�ܓ��T!�����ZnT,՘3Tn�^X�z5O��q���N���q�2;��&#i�:��W�F;�Xcsj
̆G!�htt�W픓O�o�\<M�15�T����l)�t4�R�#
pX�q�xzYM���qtt˂%v�m�]p�X	nW��"��D�4������Q��(S~d���Ș���_����G-�"�놵�0z�@H�j-���ǃ9j�H*�$R�o�m�JA,F��42�q��a�M��T �N�W���~��1��2!��y��@ ��BT����"7������S12G�~��d�@߸{H�B�Ŧl��i�j����l�J�˔h�j1��@����x1D0�� ���iLެ�H֋�h��t�PB��唴�H������}���?q��==s=����k��]"��T�S.�[���x���yѸ/�\-����}���H8�y�fxXA�9�Ax^���R�?����2٣��ʐ��>�y)V����^a*�q��t�d�V4��?��~v�/���"Z6�iF�t�%ˣ$���g�A�j��-.Vl��e㜃T,�lN��q�-��/~�s��$�/(=��fwkVD�RR5�l�m�hzl�<\�̭���Vlj2_uB
�0SԱ�� 7���
�~~��ga>��76r�޻���~kh�Q�����d���6���Amz��?��α�	�&ё)f�K9�4���J�5S*� 5�����?��������<�(Ե1	 ��Ľ'��X�H
�s$H�j�_�Kŉ�T�!��
[c�,��b!����
��:��J���ͭ��de/4j�M#�Ѡ?�n�d�����0�,�C�ϛ�;�:hʜ9s!�}�Q�����>�B»����������.�����Ǿ=ۡ(�﹞R��		��#V��K��|"<�2phN�㧞z�ML�8f�<�	�D"%�<W�Dh�)0T�M0��>}z�b�(CNJ@�㢨��q�V��[o�ZZY�2�@*i�P�4d���v��ի?z�gtM����}����x��S�f��93g����o��1����?��K%=TZ�\�7{�쮙�R��Qbȝ��ϭ��}�%
�8��a��ܴiӵ�^����o`����ip�!�DeK��'௯��ړO>�=c�lW@/^|�Y�C~
��B�R	�Se�w�}����WŢ`���|��!�Z&�c�*�N�}��4Q6�r��Q*���)�2<��t��.�ƍJ�R�:qIC��s��`~�XI����r�	'�g��'�x"�S.�W(�����ܳ� ��;�]_y�5ȰD�JeR`0zY�jU*EV(\\�e#�:n��&��v�څ�uvN�,R��F�D�[WAX����#|��p���ťqn��C<��}��R�;�n_�$^EǪ�ڑ9��䬨kN��Z�.^����V(J����D�d�(�+x��PP����A]4�90rx�g���xH*���!tx��x��nI*�(�DYD� ��ۿ����G����#>�T�5kV��_(�H�ѭz����'G�fG����S��f��L}ٲ�0�u�ؼש�<����LZ���H�*A�w3���]��i��	F���k��
C\!x3����M
8L�G��_�zْ%�?����΂�K���2�<����&���Gׯ_/N/���耇c�,("tx��{�]�p)|���̤��q�.\��UG����s�]߼���N9�t�@f�l��_�����7�XBiHv��\:��/���]z��&��Wk���f�r��WT��):<�����u�����Ĕ�xld�a�:�G��fx������~���ל��l��F�Ҕuj��ܽO�n,�J�8��JP����pl�<��7,�S��r:$4r�Ly�d��Ht�>19�/^�ȩ*���J͓�C��;���H�.Qe���c�F85�ҁ�bFR�Ns33U����HMT��A���Iǵ%)�H�@BMN�h�fnn�è���p��6!o�3O�T)s�9����j~=���ށ��r���莿�������GG�	�H�7x���������!+��?1��v���v��D5���P�Ǣ���5
��9ȶ1쑤�辧-Z��b��rŽ�)J�#�ڎ��"!*T�̑%U���a�$d���N7Th?l
O0Mb�
�\,R�1��"A1Y	���G?��*�q��*��E�y|���0Gip�S==��ɣ	M�*�#����$�3bE����d�^x���V~d����{f�������y�x�����{�yt``�)�9:Rbd3���F=ƺ�s��ʿ���<�lh?C� �ų?`��b�d��D�z��x8�� %�q=db��k�����-��B�4��#����Ԛ�(�~]��� ��+̫��z�$��C�J�'��P���˯��ןv�Y�����Jj��Dv��y���ޅ�C����"!5��58Wr�Oo��I�9���e�$��D�pntn󇿩��w�]��`��8n����4U����?y�7����V���|��o���Moܒb����B�x ���Z����ۉzpºF��<[�q4�4��aOnjJ�" �I�<�H��|�sZ�֫U,��E\��h�w���ӟ��������خ��i�aH�6ayB�/Z���������(V�p�\|���0V{�y�I~yïqA��B�Wly�۳�c�=v�Q'�<��މ�<��ø)(��7����D��y.Q�J��P8	�!@�0�`�xUW� y�`�9��<ūfZ[	�
Z����6N���U��|(����L��	�'X�Ej�0��2L���q'����6�B&�QK�-v�������lѢ0���vww7�����lSc
���c�=�{�>ܔ4�R3>���L��-+Ru�����X�v�8�cVq$%'�O��ٸq��Q�l��m�T�p��A��k�d�x7x��g�{����v��	ɗw�<p?0����@�ʀP�T�mȨ*�6
�A%����$B�l�#y�wpڙg���B=Θ1�W��~���`��E��h�I�(lXV$�!)�S��ڍ�J)B٫uRC�F�P�,���sk�B1 �O&�Uz�fT<46>i�r�"ԪEU��2�B�@l-��6�k֬�յ�z-���Ґ�D��9H�0|(�s�s(qy,"��.�iŻʥ^�I��
�VJ��
��[H&S��]��':4<>1�LAv�p��1�OĴ��R�bT*P~�����&M; "�����n���Uf�u���W7Q�B���H%��k�-W\���>�,�P�82�[�8D�}�/^���]wuu&����&�8��]�&��(Z�o�>�'�5�AVI��Уa��\��%��/X�t�h0	��� HÔhK,#�L�	W�s�|`�ar���h1M���-P6+�-6eZ�	w���.��"]�b���[7��6lxg` �b訣�Z>t�Dv ��uk�������R��z�j�|��J癯�xR*��Ν�cǎ={�<�ē��t��g��ڵk����#,X ��O�eF!`��E�&�>�짞�����3�g���<�jo۶�"Z�Tb�Y�.HMR�ga8��?��� ES��<W��x;fնX�K.����cW��j�!S���q0�+JŽ03���?�Q�(�x����K������5í�
��=00�����\~j˖-Ӧ��"��ih!�E-�&N?���^o��UG��J�y��4�cGV"��C��1���b1�k� /��c|-S0H݀<mˊ5d�K�ֶC�@�A7�H�ؒ�+ ��	�\���l��J�Dv;�,����ƕA�
�3��B���/Y�r&MA�i%��-X!�=6;�s:t���q|���a<mVw�|U�'�邱 �BR�1J��)�v�K��]}����ӯ�
��[�yo��Qz�����Ne���T��,�`h*{����֟n���_�2�����w�����q�����b6`K���r��$c-$�(*����B���m㴧w�䆁��+q�����eI�؛k*���2ufF>V88��c��A��Q�z�BDZ`�����ە�ב�3|���}{��V�p<�9�,>�Rd(h�2],	�@���U.��s!K���G��`��{�?������K/������A1-T˫p�-��S�F��ҠT��4�a�#�c��/^Z�8n��Y3��lpB��w����n��-�?0���3�沲��D���3�H��y,iH�������Ԗ��d�����y���+j�9��'|����A1[6��\�ո򧞥\�D.P��/��:x�r{��{�ҟ�{��'������F)�T�H�N��vjt�W8����Th�x�����0��k���09�w���L���o���Gb�ȣsVj�?y�h}�����_\��m�����;@�����{]ө|�`��S�x���$ȴ	n�.�H��yGY>��Ac�t�, ��UԊ��~�������d&�,,�(���y�f���Z�%����F�-����9�S�1��#�Ɇ�$3h>���R��N�6mݺu�L�\)�8�D�N,��u~Q�Ω�QA�_�����j�b�J%n���M�k1j�g��x�pc��ʪ䘏N��r�Z�YV����Y��OSB3ՀkG�J��d��⢀�ʅ�Tf�#�3��:�P]����8^��c�	k׮}���.����O?�3���B���d"�\�'�yA���H��H0�_}H^��HEEȊrA��H��,�$�������>�O��+�@���k"�0�������D�ċ�%�y��nv7w��c!P8�h'S�$�A1P�G�|zWeYm1h*4a�>��*i\ƫ�����	7��������y
�p� �J
Qf�J�%�1�2آT؝"؅�T⦐���I�b�k�˒y��zr�������
�5}���x�D��P>.�&�9G��4~#{ȩ���4�&�A���H�@��HE��Y	�I�/
���+�3!��4\���V�I�	�Ǌ��c�izQɦ o>G�tK���"�J�����Ew��f�Z��D��<Rw4g�Z���[�d���޽'v�gD�09>;%���A]4��xA���fpS�U�u&QwibmQ;$�k�Nn��%7G,/�M����<9��%Bi
�m&ކO�:%3{���3�-p�G�������R�R��u�z����WQB$^ʖ7ho��sT� ��ݳ;`�����߹s�U?�	�����X*�t�M�w�Pno����b���|ʱ�	��p�^9�S�YU"-[a5���d8���.���\r�^~��(%���	�ڷ���7�׽G�8��m.��A�*���g ���D��jΤ�,X܂�J5E���m�֣�=����^_�<�e��7�z�'���+�v����3�ȴe�q��~�����;o�����|n\�8�)*d!U�2఼�B��~�	Ǭ�߃�6m��-�6�:�@�`|zK[8�T-W��T8���<�ਆ��:(����J�Z����@�͠R
�d�zvy�����>��cө��\�3<P�Z�	��0�(�Z,����T�T��������?�>��S��_�e/K����(؇�d,Q�����<�7�jj�.�&����n�ù�^��x�@�G�)�t�-�O�������e]Q�T��BA"��������T"�'�����T�q��eBFd���9�\��h"=:<^ȖL��Nu5wԴ4�-oܺ�㧝z�/�u?ٔ��/������ȥd�in;����:M��..	Go���nj�r��h.��g���)qA���%f�H"[,�t��+�>:L/���p�����L�{��ME̎Op�D`p��ȮJ����)�h�Ԕ�t��ٽs��7���/�
ϑ��������mm�0�OQk�Ћ[=%Ő��­_��|�	-���SdՐT4�Σճ�Ԛ����Z8Q~]3�Yu(ߘ̐/�P���#P��)J"�%����M:�!({����fj�!AX��}�CS�	�ij���A�J7((R(쩔|ǥV���t�-��2{�t���yk֬��LuIWJG�m���6#��.�vJn��UdT��njJIGz�Dc�7�)������ʁN\�T��B����[������Ё�W�^�x!V�L$~�g͝�O�;�]�aeY,�se=iH��$vM8ḗ/�
���7�p̯��~1��ȀD,�2�wmr�y�j�T�E��Y$��x>��%�\"�y�P�\�۩&��@K���`������/q8X�Yg������u�]R����0�4� �&T��������:]�
K�L���C�b�|��2�T��
�3�f��U���D9
ĺ�ӑ�WN(b5y<��U��'� �� �<�sm--�")���A{�+������߸��`]q���#�|�Uo$��\d��O��V��;��%E��g�}���}��u�����ry,Ҍ�S�ۈ�*��X��o���dvr��y�]x�3k�a���MR�.a!*���ᛶ�u��l�4�<�hU��Z;/^���a�7CV"�Y�|9���!&�q���{��Z���a�b�xʅ�v��V�;���~���[o�
N���Hx�=CW��{�:cP}���lurh]Ǘ�Z�q�Ν<�Ы�!8�t:>>	�\q�
ʸT�\njx���
����fWˁN!{K��=֡�yъ�h�#b�q睦e�\����� �9��s�/�j�f��Z�p5��;�(�fv���J�b�\EdX��%��ڀ���;�D�8�C���in��=3ay<����rR��&↶!%h��{�W.[~�lFG���HGs<LCHm�8\Q��i޼]SGʣP-���-�X�d�ze=����0u@�Ȱ�U�
�"�A؂ToTh����,�O
�L�ȳ�Vhf-���=a���zL��oW�&XA�)0[���:n��	��v	�f .WcߖXE�<�Qr����ˢ�+����j!S�P�me~=���$�T�8��=�2�bΜ9P>T�,�(��@�1�o�x���%MG�Z�_|�c���+�7���A�����4n�H����/�����ȅ��[r�6f�Pv�Q��~�m��q�#���Wx?�Ž��se��J��7��Ճ����ކ���>nP�%j�(�W��,�;}v\M��5�{u���~P��+���/M�<��Vh��qS=;>|�I;PX�܂��F��CeD�0%���?����q�FP*\P��8����[m�4y���^OPm�'��XA�0}+�5ʃ�3HT�X:6�_gPܮ�3`�lذN��l�(v�Ծsr�"UÀ�����
ùN��6�����k�������Gy��s��?�p,N���L��'�*x;�Z�*5�-�%��𿐿#��M��~H�H8��b"	�U*�}� d�(R%�/�0f��K�
�?d��cr�6]-�����+�
H�m�4I�'^���[>7���J�<� 7=9�%��X%��ypN�R昋����%%h�T�u��S���L�xO� ��r������{}ݺ��o����zȀrP��ܱsgG'U��ݻ���O|"�	Of�q�:��(53X��!���IB��6#�����;��Y�͛6myq�뺡d)�`��_|١���T��B�u��	>�����`ЀO@�99n;p��Ѥ�f�l�{N҇���A$1O�i�T=��Z�	��Ql��S` �[`ߞ}8��Y3�s�W�k׮R���e�#�h�X���ţ]M�힝�c���-�!'�V���[/^0�n��72����qfKkg���@U-lZU��J�E��42�"�5�4�i�o�6SPz.g��j��W��dq��FGG4S-�k�믽�C8��G��c̚3{2;��˕F���*4V.?x>����+?�j�J�fr�0D��>����^[�6��c�կn��}��e��?��Ï>�w���y
|��K�T�RUi����"Fc!��E���L����f��l�k$<�{���B��"#ܵ��6"0���˜�ũ��Q�O�����$F��P ς�N��5-�[����qk��Ή�ὉX����)e�
�i��󄦲VO��n���M������Y,R�s�B5�
+ƓN:��SOuFO����h|��<0��۷K-���,ttB�+ſ�uJ� ����������s�R�Q�j�>���I|��d�f*Ga�$�Ty�@�OZ
w Bv�t*U���
���1�<jժ��V�7�������?�L��L<�=�	�]T�@S^�=nڹYl�*�m���F��
�� �Ղ�o#���X"M��rE�9����Z����qkX04��o�A�v������񄌶�:GR>&if�}'�ޣ@���
 :��1�@4v���gی�CX:W�(d%�
�O<ql�0��k~�K,i��༹�x��Ͽ�p��e���ؒ�Q=��2 ��ZZ��1Ȳe�J�r�!M`}�+_��w׮/\t��YA0b_\\�K�2�^�@2���
rٯ��)n?_��.��|��O�]K�C������C�:=C�>���81S	:�CC�p�_���x�=�����Ѷ�K��������,���\!LXZ~<+��`7�4I�?	*�X�)-�me�]����KV���(J~�(,.X��#I3�*�c%iP��ж�e�����퓓�O�J4�`JG)��;���СC�t�
���?8k�2��u�:���\�LM�d�!U�Ai�G�ͱb��nK�tJ�+���)��TL���4��0-��щqۭY�&�9Anrj�������hiƇ���_�t�Ma��A�5R5�#���Ǚ_�P�xd����X�*�~�6�u�x��N��nɦ�@�
K�D����N���׫
�*�ˌ���p�uu�ů���?��_�V|衇�p���ԙNl	p���LH�(���3-�]�Pa:<���	S,��R�S�sqt
�H3�0v>7�T����+ǅ�(:x� f�.�K�w1��128���s9{���H\F��]}��vL#|���>��[;�g̚��,�� ,�۵�4�\otd���B!���b�D%_-J��H���z��m꩟��f[�jo���ܣC����.I��FdP gtu��P�71�[��z2��Őθ�����\�@	w��B_p�G��c'��cǎ�;wn޼��7ޘ9wnK:M� �$7����NκZ�m��;}�gk��d��$@ 	�HQ������r	`A@.`C�"�wUzH�4R7}S���3o��9�̌�o��2;�ο���ʮ
Gch��l���qMd) �ǭ �H��N�œ2J�]#'TX�I�J8W�a�^�l���i��v��А�z�J���;M���w���D���չw��Q%�$�I�j��"dm�ũ��
Rb�R���,���j���t<����Ɠ_�@���qȂ�
5|��Ȃ�"e�Z*.� pb��O*	zb
���T�M�e�ˤ�l�R�\�6�j#n@�<�b<��*�2jdF��D��f���C�!Nn����;6�]w����4�E����6�F%ȦU,��e
P�BA�&��[�N�.p���^���\�v��l��g�-�)�����K��n�O>-�Ӆea�p�CvT�L����'O��O(��{�:s%�8�ʃ �����$ ����R:D0�JZ͐�S&h$"�AT�S&�_�3�Yq�m۶�m�H�;．���!�a�X�CCFUU5�Ɠ��3.��~q��(Ʊo�O<��o~k�ܹUQ���/|��{���9z�g���#�l߾���19�Uc� W���`��S�p�ho<��,��jkk.����*`= �(�y<�b׎ T"�Wh�V��P29���('�Q0 ����	�Ӌ/ƴ�=gFU-ա/=~%no�&0���w���bh$��Ӊ�K�r�*�X�eSIH��!B:�����%�+����<8H�R�IX1��zz��R!GI--m����H�pI�	�ۧ��r.E:�J+j�94|�n;e�rӧ�~vjG��a�IC��c�-����H�4��[�v(���Iwʔ)��&��|��Y����G��T��	�P
R�3����yH�/���c	�g�r38�.�� .��"� �|�2 �`^���k�˓յU�>뜳���[o����B���-�Rn�V�W�*��K	=��(��u��A����\K�;ա�[>m�T����z�2cz�� ����>��ǎ�o/������[[�8X�_�旸Z�Hg2�/��8}��a�ع�v>��R/��UUWc6�0L�c(��~���/e��q�U�H�H����F<������Pח����O>���q��b.f\���ۅ�~��W_��̾�������I'N�&��5!E�!P>a�r �Ω===��T�@Tғ�����x��C7NnkZn�ςS�馛~����<��k��jƴiv.����7mݺW�;��α�^x��5U1�f�jDƈ,qُ+�+��!��d�E�OfK�$ŬY�v��;802g���퐯/�N)���zI��`8L�*���BN����ag!k q��[�nݪ3Wዾ�_��F26��_� ��On\�z�1�{�u׽��[�e���o=�r$�H�<���w��d�UԶnt"Az����u�Ҋ�m!�ioo���z��MP��Ӧb^c��X�����R<FU�t��k��v�b �!�hx�
��]�܋E�[T���"�b�y睽���P-Zt������;Y*�eէ�����c�%:"�J��5��S*~Q_�yĩ�S��i��V��Q<�]%�|��cD/I��$������gN�'f��G�	�r��ݧ4�L�7�ޣk%�Y��_��c�|H$�+٤�0u�4ir<
�brת��C�~��k~�_,�>�G������'MC]�bŜ�3���� ���4�%(l=0(�j�������O�8�� ykB��T ,�����6�F[[����q�m���UB���ǯX����?��S�;[['�v����y#�wxku�`���[p�W}�s~�>䜟����A�)Y�,;��5Ԃ[(横x�E�V�ad����S���A0-���c�P��������;���˲p��eU,�� pR�	�	E�j�s�p��wjժU�ϝ8�p�B^�<�;u%
��Fc����
ZFScS"��sRѪ�}�`AGFG�zF�·�B�A6^.+~|��4�vsH-�nIzYH]�7�A���T����B1��y@8��?ۏ_ ��^��&}'G�}2:^�q�(reG\�@�y���p1�P��O�X*���s�ꈠ�OE�b�bF���?��O�(�ۏ��̔ǳ PmhTA�P��6�Y6�CQ�~�VsE"=�Z0�ݻ�R㹎�v)�P�%��lZ���Z����u|�����H(����1Z�@����nVW�_�9�q�bUՐ7�_׾}�.]z٬�k׮ݹeV��ϒB��� ���*S�`��(=��L< 5�#7/�IL�O*�B�ў�\t�W��ў�x�P�Q缆��g�n�#�Ն��o\{]8��\�����`=�3!���[nYrܢ�6�>D��oB�����1�Xu*��|��~���t9u�
z��[oݿ?�>F���/����������sO:�x4,~�SO=��7^7�r�S�L�2�S�dD�e�=��d3|r�n�sy'�@}��g�O����c�vq���B�����Hİ�_��:E�*_���3f̀V��%ƕ�Q�)l��R�<p�޽X�鬮�U	Uc�lZ���/bSg�Y���P��
��lv�t
%ϥ������87��vp-�+I}��mّ��%�&�C�p���D�"�'�4n>�*�%�$9�zQA]���S����_x� Z)�Q�'�H�]�.����쀀҉�?��+N>#�Z�fM����lAI���#AN���5�ٍS�}~\n��I^�[�ɹ�0�/���1���K.�䏿{;���Lg�JƏ(qe��*aᒑ�mO)J�	M�#��<G�eej'5���e�-]���o|]bcħ��'o��V�ZJ�ΐg�u�F�A�sR����?�U��ۀ�p]���3e��o����|P��UA�/�1v���Ǣ��.�죏>ڼi�� 
��rcM��	˗�s�9�v�"��m޼yj9pqn��8�{��k�M	;��r��SO]���o�O���	�<��Qތr�=� �jV�ܹ����$�=���S�'4�:�wހ�e�#8�x��l1ҥ��l 004��z�`���0��KD}�AQqI�d�Y����l���S�OU`�����⼐x����=D^"��r��;71�g�oK���X���ip�^Q+���Z�Z��?^��F�6S�B�RY���+j�.�6 ��	��[n�Y-Rdyhx�S��S�e�/£:wJQ�PmI^�*���cc#V����9�g.��,�-� 	���R���)H�/ ��g��1���gD+s^ţQ��w��c�:�wN����/�ӌ͢��`{�Ӻ�dGPT���^n"M\A$T'_(�R[�U��6D �(�ݼy��?@m(7��\�P3�t�l��&���!�`�B�={�����qX"��E�ܔ����p��t��w\�:����4g�T��:�����	�&	a<��I�_|ѷ��-���r�4v��?!�΅����o.�)��q�q�w��wp����O<�̍x����Q)6n��u=��e@æ��������J���	X�x���h[�ei$x0��˗���3zz���2��H�d�7�X�?�Y*B��wU���>��e�\�����z*1�|�9N ��>i�栔���,�t��1k�3����39�����{g��.�H�!� �C3g�$�px'���ϱ�.���͜<S��y��K�{�s.�*P������9�O>�w�<�0����0k�+�!d2����ݻgL�jh��r��� 3构vQ��
W6�C�@_���)����\I������hA�(s��*�l.�E�[ȣ�g�yd�dJ55�[���u말�U��b#mTk?44�.A���dɢ��*�TE���
c�h��C����+(R&j����R5�W�S�Em�i	���}�nyK-�ģ(Ƴ�K���E�L$jjk���
QT-���E|�Ĕ���-�݄�+g�r�tMJX��P�����N��1頄?��T���#TV���Ƕ�@�����L6�j�J`A@���Vp/�E�ڳkWs[�� 
�$��q��Y�a{p�,�eZ8�s��]�x�u���3r�iY�q�)�
	O��d)'�*ֵk��)�P����d2U]E�Ō���͟SUs�B0@xZq�K����_~�W��8����e�R��̎���N��*���of�W=��;ݕS�GD�eHf!�5�w�#�<�A!(��i0��몰��4WĻ�Ph���+?9]��S¼Х��7S(�PYQ~�/>��ַ�z���VzB`���tb2�w�yk���$�L2v����ڌ��(!躥R&�~I��;�'�7n��կ}XS]c�5=��sBp)V�PM(�E�|�*N��5���{O��D�(V�i�%io)&���#bkk{<^������X	�%>��d]�~�����}G`��I��qy^j1��;���פC�$|�(E}���IH�"�*9�,�%�)�Z>�w�)%�_�RG4Ӈ�Q�\�|>iRD$&	�L�H�)/S�y�Ԙ
�Zq�j��j���)���!�`4��f�?���F��U�X��_=�Ѯ}������h�!�+��B0�9cN4R�9>6��C�V�M�<��O���=��H�?e�GB�A<N�I�<�
hq��U�	)��-8�� �m��@��;;�2��0�"�h??Ws7���ڵ���:�j�3#)$��|�s����Xi���|Jϧ�[�zE!��*y$�h����X��*�K�#�(�
�kj�F������<X�A�!�ʑ#c��w_ `H�@�'�N	MmST�[M��d�7�|��1�ͅ^HY����s��F q��a#{��~bt�'[���`����)�e��Iru���I�L�fR��L$�69K�<�b���G�na���0��B�\V� ��r/�+�3%�!���W���XXq�&%�zP�C��.ԀixX����]�Y�� ��g� 9i�P�MP�֢(���sp�(�u���p����t<�V���0a��jJκ�E��RY��$�YHE�sb�򙰌�Ph�*T��V�Q)����$�� K<�z�Y!+P���.�k�e��/i�������~��#  h��a\p�?��q���ꫝ��O?�t4F�-3����e�$�Q�J��
7 �]�-ъ� ��H�a�L1�@>E�t�ѣ���L�I�p���hztb���m��h��~5*���x:;c�ȰCݽ�����oͧS��	㱱*D�
�q����̔�S5�o���νrl/ ��;�h������h���aM�5�n]���1����@_��n�T�)�9׭�
�E����]�	�;�Eʎ;������{��Y����S��
Y[hv�҇m-S�{�"�h� @�Nd�R99�u��'iW�q���O�7���V`dhD�E���,>�H�+^���i�i��#8�C����)3gN�~o���Dr0䯁������ {ry;:���=�� �5��A7>��Wҹl*�4H�D�0)�[��DZ�H�~��Ʊ�l�H4X[WEΰ|^�ȐV�����l������{�д��ӟ>ݺub4��
�.
�x���M�v���
�j�+i��}�m���)I�7�Tݒ-x0�-�_�&��CE-��`uMص͢3;�χ�$�U�)��)��}�������Q�5�EQ��@�E�U�e`D:J���B�BW� Ca�xP����:|l�HO��{;�2$�ds�p�h�L�1���������Ԝٳ!��o�Z~�����5?\C�9\�+Ln�Q�~���N�t�Zz��$r)ep����C>�{��\�21�vtLr�	l�b�͠�,+j�&�w��6������ptph���3�`p��D���X�~��w%ȃ�!\@w�qǌ��W\qEm5e�m��)��L�W�X�i�&�GR��|�	Ԁ��!I�1a;Q��Bv��CS�&�f@�2'<��?l��]��~#�ܹs��#4�����+����~[{�p{3�M;]23���3�1��mQ�"�ZMM��e��>��ª�
퍫h�R&*�G��.�O�����+����~�t�<|�~p�>8sZ�<{���[P�G�U<���W�#^U
�M���W�$4��䎹���q�Jp%(����{�����y��_�z��'� )��H�G�.UԘvF2:<&�I�
C7I�2�w�p��h�,�łt�"�����DV��;:: ��	���=�1�ܖ��<U>K�"�k�)L�:5��>�'�T n0X)���hX:�p�<�)��bw�*ť0);��rKcL�	@���^�3�M�F�����{�����0�۾�CbK`f	L�/�l۶�ȃ���*[�l�Y�9s��Ɓ����$,&e�
`��xT|&��X�9�?X�}���AX�^xKS_GHlߞ���Y���3������u���ǐNQ�l*�r��%��3|��۷͟? ���Ń���E�`��-�3�e��W����tO:��)��K�1��1&S��z衇���mӦ%��Ɏ%Ƿ[UB����������z{��Z%��6��D�r��8�ܷU-yF�F�E�%nl��6Yi�-\������`?'@��D1]}��w.��,
E�e!o�j,�$E�E��۶mkinhn��;!\(���X	!�k��{%�X�L�E%��6'$��3��~J�H>"�}�#ÿ�p�+�2�2���R�����(N�':̑a��g����#��W�V|��IE7�*�I�N��TX~�0����ٱ��y2�l���9b�p(
������ЈMI���-�m�ў>N�#���aa��������T�j!+�Ԃw�~�q�S��YNH���A5a�,O�=V�`ci$$�W��7�o�6���֜��v��z��w�>�q
DMw���7̛7o��y�t��L�9sf}��{�>܎�47ս��ښ�>G�Cs����n�Q�b(��Ed?&���r晧�p���(74"vl�rӠ�p���C8���/oݺ��k����G�c���ipJ'���k������yq���s��������J�T��.�5).	ͱ���^��)�$�L�3c8��|n�)X�Drl�dc�F"��A�M�Lqm��r����bB�PkՖv�$,R�*��dI��^����a��g�| ��\&�g����D�1�TY��=)����nĭ�Q��w���'��|�:7pf��{�b�O���ݩ8��o�:�h*FHy�c�+��-)�"���#!^��xR�Z$�Ht�T����������N1�M�7�{�RV�s�'�͘fr��� ˖-� ߰aC����f� ,3V�B��dk56F�kYal��^�M�9o~��ݣ�G�ė�5�"����BM\b�3HE;EGt5E�]�k�:n��^q��-��)D����5���N��z��,����bu-�V���iG�Dj㺲i� �[����[g�,jTU����/BC̞=�.��vX�d�?��'"��SZ��y�f(�X�����$GG|S������l�⥆O���b1꒜OR/��v 6�$U�~/�\sݤ�zHǡ������u��C@�y'��g�Ѱ����_#!5>���޽���U��(���q'tϳ)��`�9��K��;�M�8�I�Ϲ�8y��AU���CܱO׻',Yz���������?��R\ӠL��h�;3)j�J��l�����K�tr�aF��x���O<�{��L�<�~���s�����q4w�?p���qک�PF2Is�_|��G53d�N����(��	��+�s��QF���㥗hcj@8�	j9�srQ+��� ����Sy�����2��s9"^Q��:�������X��N�I�m�+&�)OE:��Sj���i_��b��s�Ν�,ot�CbF�)��}���t� Ծq&�P�C�P���y6�2{�n�\�P�*��Eo+~�����H&)�!�IwtL�oJ��}��Y��e���Q�55�Hlxt���NS�H$�h�qR%�L�l�9�2�~r�[,�C���o�Q82�b0I��b(���V�Y��t9�Xz$�=oɵ�ah�l�:�?����͛3g������-��X;:6-<��dp�5=�x	���_ex$��y|��ԋBġ�B������+�;�<�W�.�����R�,c����ȅ^�K<{�JY���$�W���W��ܳ��~;^i�ox�ר��g����#���.��X2���=j�	]��Ȳ"�*��@Bc�[+��矇�Y�|�	��CL���1��N�ZZ�551�eQ�<�2�v4".�|�Y'LI8,�dp:.��5���dM �Kf;?�p}m=׭�Rl�������i��9z`���9� ����ZC6�TN�4-?�����S�]��r�2���Y��7O�R�4���؍�+�>��T0��
�D�{e����+E�^�~�FM��3T`M��#���駟�ݽ:_*N0;����X��ο���f�cX���S%5�����ͷ�TW}���u!�vN����F�L�Ί+:g�mj��J*$$k&����;&O���׃+�V�������A�c"�kP����0�5w�/B�9rdނ������d�״����VX��(9�J9��r�r�tAg��Ef����T�������p�~`s�����֍�Z�re_�fK(^�~=5�3��e�1M���k�jZ�� 3�E���:,�\&Q��?�����;��s'M���a�a*~Ӓ��#�<
�h�ޝ8��P�9Aj+j[{;{b�g���G?�Ӥ�ayU�̛W]U��f�z�o~���3�����j�@��v�%,'H�V'Our�aqqjI����_�z���<}�)�Lni��2���˓E�;�{��X[1FX�SY�����H�
b�+̯C��.��?>����~�M�l�s6�@lٲBk��V��?���G����ItR��HL44�:�jim�#��pװ7���@b>ŝE�sN<�A\��۷o7"D��j%< bب�2�?rE+G���U�N�J}�K9����g�Z����w\�EN̤�L���	��T��W{�����򗿬X>��_�}j�(��D
���W����v͚5�����^�$���� ��٧�"
��Q���c�}%������._ �r̢�����(����:�k��Zy6_LW�������6�`ѥ,:j���#�K/����n��u�]� �P�a
�'�-��&;2�]�n���N��J7J�nų�2��,�@q�B��i�)r]N�ۄ������H��y"�N9eU~+�ش��-nQщ>��|������6�z�����p�^�\ɜ���y���z�p7�:w�LH�����L�l7��\W[�t�R�0Dz�Pɧ��ׇ%�z��/�첟��'���7��O��J���ᮮ.:��^#ݢ���D�Z֙,�[�r�(����Y�d�H�a� �cǎ/}�K6g?BAf��x)`^�\E�\2˚� ��Mn���4� V0�(�A�l�^�j��g�mORvbu=����?P�J�	�p��.`�S���퓧`e�ץɎ#��tO(�T�z&G�b�_|quU�HS�����ltKL-b*W.�Z��(�0� ��/hܨ�l���fMXq�H���"��Q�I����|��ں~?0��'��oiU22<�p ���O�n-������ޣG�2���߈;	-��d}�%9�gM�c���|�j媪𞖖\�n�aRm6wj�������;�q�ƶ�)��V.�R�h�{�+&���޵���L�S�v]ƫ��#�����SO=%%5��Rr�e0�r)=W�R�U��(�=:Z[S#|�U��R�h<�Ï���_����ajB:\U�dr{�}
-���^�,��4VX�����?��ɮ��qf���-:>>
���w�&���N���t��+8�?΍i�J��<�[r��`Ъ��?���?����m8�G�a�Te�8S K"N\-���4�;�L>��I�	�]	c���� �JR�_y�l�n���\��8���9���_ш��ka
in��9���R���/�gԴ��{�inn jC5����=�Z��wtt`���=,��Ι��［���>���?�`nh�$C�X&���?�����K.�N~��[[[)N�K�S�<�I`s0��R#�t¢6��M�t9���/����p]�W*��s҉Zb���>U[|3T�')�����c˖-�7b��8��Bؐ��ˤ&�(�O��陿�_����{�����.�=x��ӓ�C^|�)�㆚*<Rd,�_��h,82<:}Z[cS��k��k��
9- ��Q��b������&����w�T�n۱C��ք��V� �A�E#��>�����g��q\�j@p�>�H�N��dr��i"��p��	d���|�4J?��Dx��L8|�3���b��0al�L�|��Q�Boo�;�$�!�)����A5NUC�nn�bQ�v�?<�c��F��<%��t�Xj�9٘���$	����|��D���������[�Yr≸��7o�3�3�r+l��ɉ��"��i�UP٦W�&"�[R��&�к��ꫫ>��y���ԟ(�������B�O�_5�az5"NO�*�H�C���]�b&�}�r$/{��]��)B�`�����XF�`(�E���<�-�׿����-��P������E�b�s���h�[��/��Yq��B��Y�
E'�\�\"/-��*g]Wb��sF!A���t.��_ָ�������?�Lt��khj��5�\,Jg�"����W_M]�Lbj���'{�oɒ%xyRm�q��S��o��yӺ�3��;���)5�L9TL	��K���}��y�A",$���(D��,����u�`a�:��p������p�(CtT�wK�Ғz
)F8�"��[4�}U�B)�W����{Y�aʸ�bڦ�~��߿�����U�]�;EXXgp�@0���S,r�h�	I-L�1��swb�г�< \C�x<608�r�'3A9�P��Ґ��H��7"�Z?ۻܚKWQUB�t͊�O�w���^WJ���N>�wA�ܹ��~��Cs�:uuUM-ąC�ɦ�x�znU�d�n��0�P&j��8b����S�%�B�B&{t�A���h)k�Q����"�x���=��R��TW��r�[�8 юᵵ�P&3o�E�w��3�^����B&\b�J`#IU�1�L�e��l�A���uep[OE�qR2=�O���,z��~��J�
�����؞�-�=)z�"��J���|�IUoll���%L�+/n <�&�������q7GIm�O_��+�����C�0��/~E��C��ks�O��0�o~��L ,�˥L���n�y�q�
yop�����	X��j"Y��/��j�9�1��-v�Z��ڵ ���C~��l)��8AͪL��p|p���}��C�G�$ZXYp���X�J��	�ܦV؜�D
�t���s����P����4u���v����p{&��[�����/��s<�)���!?���*�Q�����-ѓP��S�vNP�E$"D �C̒&Hh3��g2�ʹ�4�����U�.�Bd�5#U�h��$y��R+�`�<�c���m�$N�����	�,����W� ~�(4aۼAK�$�l(���A�[G�Fu�K\x� ���B�����aY�(YO�y����JAh`��̳�聶��`��e��
 �@��s*Z��BB5�j�y#�� �B>���F2(Ϛ���r3�U(}���R-9��}N<@����l�]_;-J;%�#��9�OI!��u��.���뻻���h4t뭷�y�T[�#٤uU��m�ˤ%Qh.��F��a���'ONƥ�����OiX����_S�M��0�z3E�EW4� �L#��r	�̮���̈�\yXrwA�ѕ�\9�d p�I�����&�	/I��v���������Q=�\0�fȁ��qQ��w%9X2WpmY��t.��>��eE5f�8�'�����P(�L$(!�V�N-�o��Eb��K�Q))'M�]A��\�n9Ӥ�ML����F\nr�JPQ�*A�G��t�5VӇ��-�xA4��������7y�:,��^��@T��7L����r#Q]���m
�7{�1�a�Ml|ͦGF�����}����Ǝ|��_�7�ֲ��\N��?��w�RҶ�?���A+Yn���� �N��(�s�@Tr\�E��ƴ�S�rVڔ��i�TQ��Yٿk�W\q��_s�5���8Љt����T3��F�a[C�-XpLSݖ��:�3	�E��CG��̝;oN��/~񋖏���{�@��N�G�l�
E�aeѱ־�Ѵ��(|�N`�V%^Ǵ�d�BL���+S[,ӂ�	X&���6a<R`��e9T��!3J�d�r�((��(�ݔM�
���]�;�&�匟=�8X���
�U|��>u�H���܆���k��E���%녂�.�{�"&�b�_��D�I#��R6�p�1�,%s�a*Iɓ^Q*�\V2� %��Ǭ_)�XN���sv��8J�i�����UY9���_TK^\�Tm�p)��!����&�ᅎ�D�Iz��S������`�Y4�����MN��T�jƆ�L9.��T*3Y��רϠ\�����ER}��R8���*������(a��*�T<vb��s�ɢԍ���,3����9�:$$��RO�TqI���UZa���r~�\H�%(�;�ȷ��Uv��f�vR�:d`�r�i�.�V�	$����B������x��Oi�hk�7n�ɂ�M~�m���x�-[N<f.��Ų���M@���G�&jj��4ʕ��v����~�t���H���~��"��&'>�Z�.�B��	Uc`�t���/�QP �
��Y�A"�q,G�H�*��#"�JNrf���[�+�lnSW�iD=�V7ތ��ܪD������(XV�
���%�Gp�td��Gz�I�*�����@0	p���=D7:�����ޚ�{�Ṧ�=
e�p������.5- b2(�%׬8$�LFm�����9��C����Ю]]�킴�Ʉ+�~8.�`5N_�����]�w�@6�GU�lvxx%��H�4�cI��M�O���1���~���lRp\cc}U�
�g@嗊��S�S�,_�3�N��3�VJkԩ�^���q)/`���p ai&��X��� JB�c�I�=��ɥ�I��m���5�zEQ� ���O����3Q̦��5���  O8a�p�1�����$?��yԍl_��?���w^��)dRA0�]J`��N��O����M���%k'Oiim:rxT�|���S�N	��������+�P$��5=�2�$B�u��
`�Z�O��ނ��3$z�t�.L��c!<�����x!���S�PӨq. SZ��
F��*s�X�Q	�e�J��f��&҃b����Q���*��P�"���ڧ�J)F4���ĸCy�
J�*����(#��	�B�D+}*�_�hˬÜ���o�|������xTj�\t ��a3iC)�F�3`]%�Q�*�A�')� M	[qj"e�jEC�t`e�8�!�t!J�2�Pn޼��c��袋vn߈�F�x~�ۇ��$ *��L4�R�yPy{*�sQ���E-k������і�(�������:m����)SZZZ��K5u>��[k��x�ϧHռ���HMer�,�>�&�d��-5+.Qk��dl�1�t J�h�8#�"`�e���*Fc��&b�|�	!*�� ��D��rH�l)�դ2EH�2�h��4M~�����>�`����*5j�U�t^:.�2��a�`�����j�Ț`�qKݱ��*rP�bH���8�yȎ����+ʺu�۝K���{Xzl�\�ϱ�#T��LK�]ԠS����\���*>�J�F)w��g���$��-,l��t�By �ݚnҀ�Hc�Ȓwҙ0')8A5��d�sKJ��Q@\3�+�ϞֹIf��f3�znu�:C0��xز�lr|p<9��v��j9H�Su v]���s�v���m�ge�5�Ȑvu�kk�ɋӜ��%.�X�Lشgs�:@���
Uo�O��-CW��Ƭ�S�=w�
gbVuuqܺ�},_�(�To�KY��4�����ZTל�B�xS��l��FBN����E�N<n1��N��[:��[�t�4�Q����`z|֬Yo�s�7����{��BR{�t�ܮ��M�"��(��RS1|�|!��T-�RP&K��d Q%%:\]C`8��`��˜���x}>�䒔�1pt փO1p��6o�����Q�Xק%)��L'����5U�����8NR�`����&���=���H�lH�R0��յ��w&��*.dw�hz�&�H�hS��/h��p����:6w�$h�w'�4�*A$�P�s#��D�׵*P7p85�{���jl�P[��
�4_u2���0�E��-��9y��m�hß�������N:	������ڴiW��y
�N[a�ȡ���n��%Q��`��3Tۥ�h���:y��}9��Cu���\��ʽ���@�׮t��k���mw�zT�˛N�4����^��7�P�����ڪ�$̨eMM8n*PS�3�^hhkqt��������߭��D���[��Pjj�r���S9u]�#��IL�N��I�.~[M҂�mk�D��+6�p
���B�K�f}Z�=����|f%�N��8���ofSy�~�o۶M�V^x�E��Nd)7@����g�ˑt��|�x<1:
��׿�u���@�;w�ļ��R���Q<�(���Û7o��š.:D�F+yE���=���P!����Ea�޽Lg�Rz@(��ɉq���#���������*^q���OK�G������Wݾc�����S�QR5�ᑃ����Aی��6L��8}��CG���{���{�n���-�u��Z�C%�UQK�pPJx��Q�;����0����k��&ͣS%Z8H�~�OGb1�R�Ԁ�I"Ykk���;[�)S�����P���^{-������w����h�q,��r�IQ߻W��S�Ә����#�E��{��@�[��4/�9��?�&�"���'�����b��Y�ִ�?g�vQ �TBQX�
���9���#�ݳg�9��v�abyBMͭD7��k4@��O��h�
�>LS�	���eɩ�. Fg �)�R�".���4*�{�u)�s����n�߿ρ�� �5Nr�Uv2��-��GW݁L8��n�J�a�[BŌׯ_��K/�	����vAul�*^G_WL��������������>46�ln�<������%/�X��N+4�b��u�Y_�җ>��C^I���)1,�|���w�w��]�É'��l�	8d8s���ʢyK~�`,�����_�i��.����<���Wa�۷o��ǫ��/�˸�,�я��>�����{.�>�L�#�VC��/|��Eㄺ�g���O;�4hs��tG�F}�U��ͦ_WԖƦb�
&���P�a��?��;:�g[xth��q��=$��PH�ع\>�J%g����!Bt��P�`��~{��7m����J[�������{���榓)�z(x6D8_��G�5a��w%4���}�Fa�H6G�?�ź�@�L<)�T$��ҧ�=p 言x�D8��T�B��툣� �1]�QN|�����7VSC��H��G�S�cs3.�_	�~Ȼ�lv����*%I��h	�$u\��=��_�����=Ʊ�k�믿�uێ����S�!xz�{HϨ����&���&~r;G$J>����Fc]�HJ򵄢78�,6� � �^j�GֳɍMti�ZJ�*��y�7�W^y���[qOYq&���S͇���l�{��}R�]������]���ꪯ|�+����������*��A�T�ױ������~�w���Ж*1�D�S��0f�qy$]��c4�ܧ��?�c	h�p$J�#��_���?�k|	6��`��O���˯��<���;4	&��/~V�ѣ=kn�s���O=�TM'��w֮���Ě�}ph��{����ĥ���C��y�!��[p�v�����O�*�:�����iб�R4�����Ԗ��M�0�����~�?!��q�9:�� �y�&�@bm�����+WNd�M�6�2ٙYOf_H�����,���s��q�o�]<1Be>sƌ����^ �Co�۳�<WȊ�C����G�*�-*- ����fE�̞=�S8f�����:,S|�*�p�\O�n2�[j�̙��@���=__G��\VΏT��V�X���RX�dI�:�еe����څ��k��XF��/��R�ʹa%�es,ַ���e˖�M}hx��>��~�wn��_�馛�,I�`�Q�&�q�>�^���E�P-����:����?r��s�=�λo�ų�RH�U@�J;�����4�[
|e2䙴��U�k
y��_�fc��{?&�륺���):�|�2�˸6n�T��[�9>[���pi�.�9�چ-z��vڴi{���iii���bkk[}m#����X2�?��s�p�䩳�����Q�Jս���Vҩ��05��O�ӿ�� �DC� 6�}�6����������\r	��� ��.���u�<�vz��V�>c�捐m��|p��Ş��ڱ���w����3O�w�yܳ��=�-Zh�i�F��~��BTBH�yWW���ߘ�f����@4���Ga>1���'�G����_m�$kM�����u�|K�MX�ϟu�`_4jf2i,��7��'@@�|�"��.�z����?�1�uh�?���S.���̀�p2����/|�L�]��J�ǧ�?k���f����7����9�����""�@(��c���Q>۱�2r]%.%:��	�� q
�E�!<V;~���C4�-c˖�W]�u�0	��$����4���+���+ =D򆃾x4���N�^~��?��O�={ �,͊E��_�l�d"I,�LK��6�����w��AlFsC='�2@)��S?�r��s��%$P2��nڰ��K/���_�\\`Re�=pB�������˔��5lT�JՃ.�H���+x�w/��
����b��]�cw�}7��B����p0b͜� �8���B�R�P��/�SH�G)SG�[��=�����g��΅jfv΄����؏�{ɉ7<����o���J���i��J�C������05�J�6�g�`!����s �ن����[x���%=7�mٲ�1<4�>u*N���~���A���47�d�}���Ã�5�z�К5��SO=�3{�	Y�Ѐo�}x��1����w��ð��G}tμ���P_/�B�(��� �X�q%&��VUdq�(v�S^�^�D~���r�)c�}���g++���l�4	����q���Ǹy���!J�	���S1�=��&j��6��g6N�0�O&n���f�֦�e�L�`K���S�0���{��IKdDy�G�b_ �k���o�ᡇ<�s{?\�;��,\����?���V�:��#)�������6Ò�t�IX�O>�rJ,{�&���	Ca��Q���o$V+�gňD����o�����[o��޽o/,�-7�N�h��}&��Cc`2	�4���􏏍ێ2gΜMB�5��#�1���U322�$~�R�ɢ�pQRI�g)g������a��.jDԋ��J�p�
���j�j��%D�Q`x���Mj�4>��L#���\C�a��I�⾾>|�H�~�Y~1�8��͛И�/�M�2ɬ�~]��=�3��$���[��a�x��U*2��d�R�m� �FpK	X&��ȥ��<��S<�&�T�Ν�������G��,v"�=g��<�"e��OHu�ή�uW8�2�����0:1~�]wI��@	CKC��~���%�+u��N��� V!Ꝩ��/�,���v���5t͜5�/��7�X���Hm	��������DM��E@��L
�t_ׁ����������>���2��5�N��駪I}ŦdA�1�EP��)���<7o#aaY��*n#MB�%���u����@T�����0_�r�:��|�ed�J~J�^ �Md������Ɔ�o��O?!x�5W~���}��W�����qrk��n�k��;�SyG0�����oۼ~�ܹ�F��p����}��f��=��\�����	8ܸQ@�'�|2��w�{_��dq�q٨�&_��0��������+.{����%ĊL�T:66}���J���,1����=v�:E��Z��Ʒ�Ҹ�/^QY�G_f��<$�I(0V��5�$�N	�n���犀�3;͝;u���$U`oP��Qj�(�Ƹ6�7�x#�����C�)�V%;!��N�S�-[6џ8+b��Ex��!h��cn�Pj�(L$?�#�nWٸr�w�$��uR� ���]�_�jz�g���\-�f��$1,8^��a���χ���u3�j\w���8)��3e��3�<C�8#?�M�t�H����V�1W�<�϶a9�&��^Zz�q ����O���0ހ��{C=�9u5Uk֬����"8Ի��"����,���!Ad�)g��+�p��$���VJ[�il�l�2N�B��cZ@.s+�*y��Q�%�vǁr#��V"���~�`Q|�ڵkq�n����$'&e6���s`���h��V����̞=B���! �_z<l�����8�jd�����\xᅇz{�wm��.Iԑk׾�������2CD>^�.��{���1kŲ0I�@@2ӡy��{wu)>vLG����o �`�(��V
�y�4�Jȍ�n�1���i�%���FT<��O?mj��u�^�կ~5�7\�U��f�ne�N8d�D%�b��;����ħs���9:ꔆ��ㇷ]�5f��F�.�(�ύt��`�e�;�G�f�t&
���8�aтy
�P��0#P�d*��a���K"���b�J�K���s�� �N�9(�R�*1k�Kx�H�IR�XT��oM��[�SY�S��U����KS���d����Z�l.������$.3����㘛�k�#u�̚9k��� �5�W]U����鈛���ȁ�I�r��CV@�]����Bz`�ǲ���������t�b�(��D�� �R
����$DՔ��ے�������Hʡ�RY"AI��t�{l1��"~���S��T���QU@zL�.Ǣ��mrk���O��p���C!��X@�L*���Sh��_z	��k'MOnظuŊ�t�-��7m�ڹ�(����D'�j�$�~�zL }Ŋ>�bz�]���Câ��� ���o�}��	)W70��)�$�ƓO>�>��+矷x�؉w�y'¹��iGR�p��rk�W��1��P���F)q�'��vu��ǩI���[�QY�]���"
X��uQ�x���%�LiZ���D��������� �����w���Do�!q�C����	��1Y���r�x5�g��w�%�����{��͛w�فqJ"��J�^��9�u���Z�ܰ�D�k�)��j`b4���L�7�r�[`N�i )�`vR% ��:�Ik�e B$qW6Y��u�"�k�f��%;�*�I�魭-dK���T&Mrĵ�RrnqZE"�>
G"w�q�	��Pzm:�1�x-ic�6T���ɞM����-+�����L[N�?�M���W�F��K�%)L�+�.����Z0���T�T���}1|�d�ȥ�U>��O�FL�2�
�&uա�.���l��n�ԬNt����~\�W�7)���4������}��߽{�ѣ}�z8^1�%F8�:ib[cL�æ'RI�D��-��͚>_048�{'9X'5,2���a.	K����=���>��=��|��'��f�%�ɀOO\v��q۔V�3��P59:F���]�$t1�b�v����s�=���):" ������m7E��k�N�4�GLgՓ��6Ǜ`S"�,��;�fƱ8t����o��Yg�~������~��xmv�-X�r�I%M9�rk�5=��A�sg�+���#�{dÆ�}�Ū�j�X�S�T��v�*���c}X!ԩ��H�Fp�V�Jm߶�`�L�v�k��sLJ�����h6C�1�A���6�@�T&&������J�x��%���E]��k�m۶�Ȕ�mݺ��跂:�p��h$��J��}�i�aҤf���o�k�	'���}};�*��{�&���:������2����Zmh�#���x(˦uX��ɗ�[6s�@�� ,�ƈ;�:*f�9bʡ
zQ)%	�TJg#���X�gS��Yvz��;w������R���k)f3ٛ�k���of1A��o"�����G�y�Huwwwu�7w6����"d]]24�?sVg4��9Z�P���o�������hW)H^L�r��-�ƪ �}�c�L��B��$�@O�46��ia;�|W�db��TBRd� QeR�7Չ8%Lq�`�}�ݻ���z�H'���^y���v��D�Ćʁx�o�j���"�����C	a9��������@� u~785�����͘=���L"�M�&8��gg�&�A��bMI~l2�ڱcV�D��
#�q��h��x�4p�1�@�ǋ�.���vwq�0�`�B���\Jh���׸�[,��s�[�?��5'��+7I�L���TN\ǋ�LJ�%�m�$u����.d��#Z)/Y�$gx�Q^Ƕ1$X�P�l�A8���]�?�[�>��>�&��_|�ː�+\v�꺺U�V��@�{{zV�Z��/_x�'<w"A���+KZ&5Bpmⱪ�Ԃ�������4�R_:����9���*x��2U����Ju9�_+�d��1�,� �ܙ�h�г���9z�0sU,"����s2�C�J3n��裏���.�qR�&I�_�n�ysE�BLk�d��n�໲Y*�T��)\���0q��ei³JSP����8���>��ֶֆ�z�cs4�_��*Tz���J�ǖf�h(`=��ӯ��
fF��ur�!��+�+�S��;g�hD�J`�mm�C�f�ƌ�O<�dg�t&���4��۸q�/��W�z��plڮ.j���ko9�sN;c	�Y�HΛ�����`�-�g��N>��Djkj���{�׿�s���Z�L�+�5��(�bk��itsY��}��/SpM3 s���-��r��>��Ch�\K�r���8�Q,Wly*��pAm��ͪ�D7���	��B�R��E$�D�key�,�G�M��|�l��dF٩SHg�*�r]N��߳���ݻ�J^0<W�~ـK8m���~��=����uh`���n����Bel��?���w�w߽߿�0v!^���ZXk��q�UW�c��+ON�ΕW_t��z'��G�g�]�0�\���\��|Z��ȑ3�<���o@".�3�����%n^SMP߰N��Q�W ��X4���na�rz��7�ڳgP4|29��+A��W�f&XC�d,vS�N#a2mL�l"J:t���+�wo���ZDf*���L���W���
�ϴ�<��`84s֌���,���p"��	�`2q��Y�0�h$*%�;(6<L�n��k�.$i}�	8��oݺU7Ie�Um��mP���8f�O�c���C[~,��M����ꡑ���6���
K+�����\'�K��{�3fL�#ΜA�.>�� <aCe2��˗/_�n�n�����$И�,ͤ����d�Iu5����$dR�gED�P���%�a2CԞ���/����J�����׿RbgM}�\�&�˥���!fA.8&/OP�L}�$�9"s������.p@���a�128�lٲn�&�۷d��瀩��\�D6!u���a�J��u����Z~�J�[�l�wQ�&lB�R�d^����qꪘ	���ٽ���xq����b�G�v
 F%�{��m�>���T���2h��������?t���ߞ{g,V5���y��8�t�MEb|�JQ!P�z��+O^~�%�H~���`)d�e��?r[pt�4���lL�����GF��4#X�ļ���n��NZQ�L��.�.7wV�c!s�gs�x|p�rSo���G��~��a�c�հ!���}��:;;	��֢E��n����/�s�
ZL���M�dC���<ҼRf��c��O�b�o߾}�����{����?t+6~jKK0PT?�/�'�O���G�̭���i>k�?��l�<��&3C}�8��^z	d�~�{���'$�(�p�4�v�z(X�2�m�%�r�r<�mJ3���f���0�Μ}�ٿ��cbSuw�
Q���7|*]ϡ����TB��fW[+q|XI~�/
���J"o��8qΰ�рE�;a�Ҷ���j�>88|4^yʩ��>\��O8�ȡ����J%>Ϛ����,DE	�����L�6��.�Q8��e����7��V�h�AP��G���Zۊ��ۅ�@�%��zہ
w�)d� �f�7�x�e' Njnڴi�'}����
0�ʳ������H�P.��B�8EJ�"m��E
-�#�R܊�@	N� ��n�����q9gf�?�3�_��+W�̞���r?�'�����ǢxruE%��h��4����|�����
1���ʦ�$Umnj�����QK��w����g_BD���(($���:C �di8#Љ�fV`��"܇`�b��tC�i!��>��nhk���sϵ�6^y��>�E�䓗y�O��^z	,�����݉{9�����_��!{����h��[`�
�Ն�����0�a�R�&��x7@�j`&�T������VPء��ZP,9J�T�˕�k�AHx�ʕ_@I�����,��M�:��O?���e�V�qshT�%��wn�ۿ/Л�d�D\'��ݼ��;?��/��2x�3f�}b:��%~(kc��q0XwW��sK�p/�GG�n�=���u�5������y睷|�2�c�(��n'�'�	'[�x��@!�|X������{��ݺy34�)"�S��Ɲ��	ʫ.Z�"�'� ��;��:�Ϲ��c�
��n�����}�b��O?}�UW���?_��?<� h�ԏ���
�H�@�\Vo)/�HS`�9H��c��iD�a���<��_�[���d.��	$\�6.'k���Pq'!�yP��%yA��Cl)�]x\T����߿�Ξ=f�(1ɳi��	�N�c܃Q�#�J���C �R�� A\��;�a�
�z �x"%��r?]=�h�'��P���zբ8T�r	l�@���D��br#���/���ŋw�&m�͍�h�jM���ܶ�k��dsFOë�|��y�Z��:�,���'��?�"���9���h�v�%���~�	'� ����q�Xܝ3�8���-:��qq�������t����I'GF#'�xB�2ݰ���
��޼�*���ٵkٲe,.qV�F����!�R)�)?�%����𴲫W��]Y���$O������#����j�����)�vg)XG��f2~�R�RO>���O<2u��<l(��zݸ7I�;�π����o\z��Y+���'�G����w����A�Y�}$ҦFm����Uh/�:�uU7dR��-(���>���h��z]�q+��gK���Ɔ�S�.}���{z�Ξ��r�r�$3�!ڣf��� D3=s��Xl���|��O�?�i%n���`�K0G�H��h��>��ug�\�2�Ը��T	W�:X�gktp�>��&�������WWC>��+���I�$���2
'��.7�܁ q�]wݵ�{7li\���  {�硢v]s�|.�w�?��w�w��λ�|�e,�kiN�i�[#e�	�C���s���>�L���[/��*��!�2<k�s�r�N�lo����dW%8g9�JM �$!�S������ܭD��Y���$[���X$�vQ�I��* bg����0�(����rX�A�H,Se<�/2�?t�\�˂jg��ޮ�i��'{�t�|�Os��x*�܋/����Ʀp�o��-��#�w�Ԗ�~r�{o����:i��.~w���Gw�q�a�z����x㍷�z+.���_�����߸a-�[|nW��:%*�ɋK&h�.�-ʈ:�w	�Qy��'�U�
�H�az\{��5uM4���5=XV�kG�����S��H����:�&���=NU��T箽kV�6}�澱A2p=�-�fh ��س�>{饗��u4�)�V��d�Mxff��'����;���9�,�>�����8�O?�x�ҥ`����w�0E!�h�5'4Ķ�h�Bu9g渶���h&6�mn�.P��+���!i|�	����k�[��9̏SN>�W��5q���E��z�	��{�y��,�R������2@PsK�1Mb�)q�R�rn���2�%#�?"wG�Z��+�^����Sr5��E����'�8��ڵkS�$�A��6���iݺu91��q�$]�2eb�қo���ϛ7�i�ڵ�T����F�S���P�'��Cx�1(=����|F�3N��@�s�@�D�X!��Y� Dp��#��E�f,efL��,��t�T7V4i:�6+�7��TM���3�A��2Y���1F#Q��J�{�^��d�K�V}�vժi3g��/�{�5���ǜ�A���s.����>���y�]�?�|�"��/��g�������=�L�5Ǝ�I�f�x=��>Xb�\|�w/!�p����oD�%J�\����̙c|&ۦ�?��ʕ+���=�\�^(:<����"8��:3�C~���	
��)�E��p)���A�ӵ�s�K�>�䘣O<�Ă�oh�mi��^�`��7�=��{����C�9�tv�(�+��&��D�z���������˞}����Qs��=��~��"F,q��(L7���%X>2k�OE$+�� �{�z��8F���'��v�ؑN�~�����v�HWW��3]��7���۝(d�c�ᲲВ%���ڶm����߿i�֕_}�j�$��?'� �a��E�&�F4��d�����������ƿ^��k�� ��������$t�$�3(Q!l_����"	��@����UlN?�U8R���Uv&��@�S!�?��@mmm�c4~l�̙`Եk�p�h^t��p�s��`�d�`y9a(���|fҙI�@���D(��͸e�R����m����uv����)N,�&�D����8��JeJ�bdZb\�%F��R	��"x ��ӟ��>tѢ�O=uO�lOz��͜	+����_���=�,ڶe��goܸ�$]��wO������ᅂ'����9?T��ǣPd�;]��Ƣ!:����{���n���O�q��ؘ�s`���#𲝢����2�'�x����8����B�I̲ۼaͿ����ؒ��{���t�?׶�.9h�z�~hdx͚5up�46����q���#����-�M�5,���|H�}Qڲu�.p�ZQ��_��<��p^�4p2qP���c���>��` Cӹ���j>?�K�����I��?��D�;������-���C���7Ö�k)�oh&v�̃n���i�5�W_}��?l�LU_���z(M�O�`׈A<G���F�|���H�	�¶h�v�bŊ/>����� ����jƔ&@�m�ie��eύk_�#
�ETi/�U���8k�  �l��x^9�<�������`b��vP6TwZ����'����I�+�]q���l�&X��KT#RW�0"ryb��$� ^g��t2D��S4�rA"���	����U�"�cL�(���9B{CF�l���˻n��G��jժ����/��/w�E ���ѦM?�0ͨ�� �RJ�1o�Y�Cz�?���� ��Xj_�%�R��\X�iF.K���E(Շk=���wvv�W��|�W^y%��eyĭ9ƑL~����}{{{GG{SS�&���Ѿ�;w�t�p8�Hm����j�h�K�GEپ}h8\5�U �o��Y� ��Q�_���nΜ�4���˽�}��u�E����x0�7Y�}U��{��y���@�����b�4��_']�L��	��&@A4�P��ch���@fAA�b�~�/����ҫ��f��Y� �f^r{��t�c!���ah
$���#Й�� ����w^Rq�pW�R�,H�d��WU�=���t*/PL��ᑈP2�w�yoh�ohx��e�9���À��l�*y�\�':��0*Bu)�K�,�@�PU:��
��s� �:��SI��@�T������C�@6��9�̵i^�u� �iy\�t��]`T�m�M���W~�����f���ZTkN��/���I3/0������x�1�g�g �B��G�>�!�_Q2y�|��F�G�����_�$���l.�Lq��谡O;�uM�B:m���p(�chh�����^y�������<nϟo�upό��"��������̟��؟9�i%(XO&���1U3�5���|oMw;�xoA�@VA���({v"|�t��W_r��bAJ������oV��B-��T��qq�8��ʱ����z:w���;�u�R�DZ��\��v��j0xY'�S�r��UEƢl���`����H�{��S�܇��1U~�(V�P$1�X�/S��'p��=�,��)��R��8�9�b��MZD�@�&͖'�	^͜��@��w�Ǒe��i�_�^��S�!D	wi1`���D4b���j<���jf��(�27n���a��%���4)%��B���8�� �09��6�D	��ꚨ��&}I�� �S0@`J������?5�͎;��a���$$����!y5Y*�v���e�]�U���k�u.:}�zK���Pb��OP��/�\_� �}Og'�Zf���	[�]���mQ�uV���y�-�����88�I6�)ajװ���`<.(c��2.{eV^:��%6l�d�  ��7�'n�������jim���;`~6�}��w%�P:mZ��G{{<��ӡ*�뮐�Q�F#c�e�.����	D��'���F5�B��P���?[S+��X+�B�r;|mc#�2h �� ��5�A�6L�m�R�5�d���h�GT�@#�z �|��R^�R����3���"]�d������o#�o����Ͱ%�5ɰQ�C�.�u���ҬY�UU6��O p3����ry�^	�����{�9���E�D��'�ս�����P�$�˖����G�?������nO^dde�K�4�ײ��9Bs���ϟ�/oٺ�c��/ �/�)�QQ��pD�BFx>�c�ewyEճϽp��h�w��AUĻ5�*0R��[�d�Q*DN�����	���E29�!�qҙ�J�/�X\��<�@v�\���"gr���1�:�E�eF#c�,\�����g*�e�5M&�H]^�-�� ����}>����
��^�4M��cL@B
�'J_1�T	,GU&1��v�ڲ��q��̋1\��v�~&�l^�B�#�Ψ-3)2���h6��V�=��o0P�v횛n�b������F���.?���aE�?���C���m�^s�)��r�m>�à������o�}��s�@$�ׯ��_���w씶֜�����T� ��&�E���}d2A��/$R�.˶t��)ZDti�	\s�����bA��e� �[����0-���b�nUsЀ0&������y)G�h���ҩ�17�Q��Gv��!�/�H�|����Bv��s���J�y\����9h!H�9s����*��%P�IOR�����SOA�oٸa�̙{�:{�1x2��9�3�,m��E�NV&3����n���C=��SOݹc����Ǌ
j�K$�3�U-�L��;��<>��K��!b.��R8*��\������tM�*�N(��r�ԜKxG�4��8�0�Y*�E�=�'���=���(,��Wd�Z��v���]�A�}��1��ؒgq�\q�M�o�ĬR��mo����0�D\��g�=Yb�s1 ӆ�� ��5�f.?Y�ȑ9�����o��U���T��h�b}M,�k����� l��g�پ}{sS+����s�}�}����>oy뭷���_�@�lx�K�?��7ߜy�UU���>�L6%&~4��j�59u*��-�im+�N]`E+�1|��x�>�E���ɾ'���_"?1��e�o��' �5؃�����Tu�r��|p��	�&�"}��p�E��0�7pR¦��.�)�S��v0+RU{2^r &.N�d;	B(�J���pY�ko��Ti۶-������Q�]��x������SZ?��PMU�uJk����?�|
�iikM���X�Nw���T��ZN��H��h:��,9��'�~zǮ�\y�r��R*4!��ͥ3d��]�v����}��7�p��fi��$��L�ڹ�{�N�D�ͦ�<��	K��D�='�QDJжK�7q0P���+����� պC����h����3i�9f.�V$��O>��*����v���E��"�0q����(�6l�j��\��̜%"�27��@"�٢as��s���qrY֖HF	 J������L�E��Ŋ�z;�N�1�����P� 5���ѢN���߀�
^R��M������`b@����'<=Oss�*+c�Hue��0֭[���>��9�T�W��Z�n��?L�ڤ�h]8�h\�w�,8�����P���lp���2j[ �q��Z�L����s)��8�������kF�"��g�נ�𗴸n�6T�4XcB�"�N�Y���&Y�q���J�P��q�'6��͔\Ј}N�ɥs�\�¤�e�`6�.�¦�&Q��y�ܐ ��v�B��|�GST�2�����00<L��:��=�����'A�c�����e�2��rh:� I]��׮�t �Z������8��t6��\y��2��'���Yv���"�Y�*����0��`S]�1�p��组�/SdO�<�b$M�1�}t �vtt`������� (�h���p��[I��v��r?$����=�g%l3��b�]X-�A X�?�׭^-�T.�;t�a)d�D
���b=5B��G�n�e���� ��Ѝd�"���>}:�V)�e��O�&�G��/�.�~uum+j� ����1F=������I�"���N.~\8<�/�f�$ț���M�JɈ�H�Z�c�UE2��E��wg������S�c4؃ŉ1,BW�|&Ϲ#Q-��OKg2��Ca��n1��4�2o��LL-�NV��"��[{��K�^�v)j�"�B��	�
D�v��EE�4񸻻ԯLL��2���F ���J�E����r�X�a��vi�+ga�Ru�e�����>�"�#�=)H���e~�26>����Vw9="�L#_�V�[n>�������nhj�(�X�,LL�� �eY��BT#L��|�d;��Ԁ�r��uD��`IФ2�bކ�ġ���t
uc�A2"�U�*P��I�vQ슪���ILV���U����X�����"pq���'���A╊oK�3+Fa�<ҧ0)gy���]VV�v�Z+�:��>d5߈��\V�%�O���?�f ���L& ȇ�PL>�>'�A	�DL�� �_���R䑑!�.�!��VA��T00�D�u�?���O]��=����{��������2z�p��v.ڞ@#�oQ�Pޢ�.6 a#ΞT�]#QUI�P�G:S�c��j	_���#_�|o[{�-5���nbS��d����ٗ˦)�Ѓ��(�%�t(�@�d�A���W&&O�w?�d�4�4�<��{�9�K����䤈O��&�4�Hc���$x�J��X������c4Bk��VE�T�+�HqϾ����/��r��*E�H��Mš��`�]}�����ʗ�����9��U��Oȹ��I'���{Ys��fN$v�����Pkl�E�4� ��]*� �\�˂y]��,j"�Y/>I<���A19� �!?K"x&�(1|.E�=L&Ιp%�kl{ۓ��}�I���%8v*X���±lذ������8��3�Hsy]��M����t��_xᅬ�	Pg����?k$.G��9���c"dPܻwo��a_����mَmimKPŬ�\_,f˖-��!� �XЈJQ��sb4�Z��~�v�G����4�!��Q�&�U�P�K���`��t&���ǵj��i_�i�؂�|~���=iӂSl	n��S�(��i!�!�h�Q���q��YZh	�EB4�N(TƈT�I�.�g�Ku[�ޣxBf|�Q5/'4gΜ���ɾ馛`a��:Rm���WLƪ�絵��������qEYW�� RH$��$A�P���[~��_mټe���䑖�EiU��W5�-���=�Щ'��_��p[KS&M�l0l�IR&�}��MFu<�9�Gtlp��#�4��\��J'<^��A��?��~N)�L��^�KXF8�O���� �1yU$TTߦ���*�L�p9A�X����,�XAh�h"���\y"&H��Ùa�h�}:]��ȓ$��&��IE'8V���;��$�������p.\�𩧞
���?�ϭ۶�o�#xy6�E#�>��S���E��v�m��J�>D�$��O��e8��1��O>Aɳ!V��Q<�iP-A]M=�ͦ�_�j�e���|��_���e�0<�k�J�Q�/���=Ys��Knaf�*�O�d.����T�.c:2��4����L���*�*|f�`6�}�d��n
!��`J4K�[��$B(P+n6��� f��Kf
�ژ=N�C��4_�|��t�
D�PVh�L�T��QGBԧ� /�-\�B�E.M���_3
+}ή�*e�K�:������?���ʊl�<�93��o��ψ ͩ�E=עK��o�ݴi�P��4g{)�K�X�)l���oX��ꫯ��sn��{���:o��od���vd%�]w��O�ϝw�I"�^�t{9%M���aE� ���~�,tD�F5�dD��)E�L7 ��+�iV�>�J��o�r��BE�ؠX�޾�ē���8|1N��������l�+�(�i����(@��py��~��Gs9RBTE�N���}��w�埃��!�u�'MbA��̕���<��������{�G�I:ܙ���0=�����q��W��_�ڱm�娢͂�2I�/�<��ҥKE��r8��ɥ	���/e�>����v�jq���G},��z�:�l���?=?�g���;���P&��ق`K+���a;,�6o����~��������k����}Y�ĭZ���K/��u���ȾB�� 4>��[�{��KR7P-�~E:��ڽ;
+�9j���Hnln%��s�#�%�X�dR汉\;��{��E�x\�=��p���E��W`{��|͚~�p�	!�"���˛6נ��}���#;������۶m;��% e,X�\dޘ�D(���t�p5���ma���>��SpK}C=���Qn۾��t��Ð͝��w��s�����'���K�(ʪ*�� q��T��dg�xS�ۆ�!���6��-e!5AU�<K'b���k��fǎg�u�+���嗟G��$ꮔ%!ʹ�h��D�͛w�E��`�}��'/����hd$5ͧS�Ds;qM3gN��q9���w�������K��"��^z.�wy=�򢌎��yvx�0�o��R��~�H�T�h@��Ϋ4c���mwgg2Nq $2���a���쫭�������pv1�CS�����|�]�	>��A#�����T�qy!�zGE]>���pف�ӳW�u�Ё�t4L�S)0G)�"`�)
g�	,��H-���h/�1b?�;��������cx1��a��L#8PL̀����>�(E��ݸnKO6UX����N�������*fJ=�bL���������rP�{��I���V|�!$4�|i� t!�98��{ƌ� VA��!Eq�����{DM`�rc��!�T�wS,'^V���ukk+n���*�W>��36m�d�I�0ć�Yt0�0~;�4����H��J���E�&�0����G�=�{׮]x�#�<��o|���C ��*�íШb���L7^o@�Y���f��B	�����Hɣ������!����+��-�Mak�_��&i��y�3�<��`;X-V����e�ٖ�����2x��E�c��[6�i\��GQSD�y�v�H5O�1|�*A*Y'pĈ��4Q+Z�I&$�M�|�h8�\:}�P���~�>�O�W\�[�O�l���Z�t82D0���� e��(M �e��>��#<�}j�w�tڏ?����=�PD��2�����Y�_��tu�$�F����m���I�����ظ!�j��EA����:� j:�f��`�XÔ)S���8���R/K|��[��?|��K/)��t.��q�y_����`��t.o]{��]tL�l�H��pq��K:�䓺�v��x�՗uU���� �c��/X��w�:o�C��g�E�����		�(`�tU��˞��c(��]���MgQ��Nɥ�^Iw�,�dMY�qiH�	/ų�ޡ!y��V,�\y��F������
��݊ýxɱ^z��?�%[�ݠ�L���M����H4p)��Ok��;��,Ь�5w�m�����R[0���;��e��!�=�PD���rn��g��f9��b���H4��Ӕ/º��"u��fd���@*m
���-�<�`Nv�A"^Y���C��<��{_SӀ'Ey [h��S��mT�I��>�����Z��\���%�aC�j#�'\U�e|a���;��x��r�7���b  ��IDAT���l*�ԕ!��@���'�|��x����~�u��l�0riڅSv;=ΜN��K���UF�)�tÙH�i*A�rJ.#�E0:���3u��G���Q�O#��ִ/{��˼�d���	����Qn���;�|՝�����u>o ?�˔�U��ܷc��߬��Oi_�f��kkj�8�t*��"�w:���=ٌ��R�<�p�����삥*&n�H�DԱ�n�W]u-Z�2fr�g�
����X�v-�>�����06l�<{�<p��㏧���xl$2����z��k�;�vс�4�=���#���
WE17�I)�&tT������Q�r�-�_~���ذq�$�Bf�y��Ӹ�g�}����[n�9��ə�ْ�y��7U�r�;��#��p��9/%�B�/Y��Ϧ�W]8ٜ�;��=��^.����E]Ն�{��EX3�b)��Bt�hX�E�	����%Y��n層8V����x��?��J���L$/����8��S�B��QJ=S$�.�}��R���R�d{�39v���@T{��
`X�js�<$E�!��W�D}n��D�E@8���I&�tM�p�˨^�_8t�e�:J�=GJ�	a�L΢�9�NL����t2�m���2b~p�H��x<!Fܑa��Q���H�Ҹ\�P��A$����f,&3 ����i
G��9�ws�ND��F|~�4$��6��>�C(��4��GU��_���-//�kd&t��>�Oi�/B����\��/�l6��qn�819��+:�bѱc�;��,����%(f]�5���hn���sx�P�=�{<찧�z��?�@ӂ��h�	�;CCC�ہ�
(!EK���i)1Ξ�?���0s/�䒫���f�P?�i�fV��
�����/R����]����{�v9����$�D�Z��^��k+�/��-S��������#����"��h v-g�c
yТ���Oy�0:a���,��G��[�����뭯�ɤ���1�J;]�?9������*s9T��O�gs�������M&�2l'+K9;�k�v>�I�
�����|�9���)A�ۣ��֡��3R�X���͘iŪU����ȅS��p��P幞�>�3�&�;��z��4I��4 �Px���@L$�����jHi+�o��-�ۄ��f�[��K���"k2U��T%��&t'S̴x��a�RiN�C��T�����,���d*�%l�B&��˯�-<rG�IČJ
ۤ2Im�8�+:!��
9^R���s�ZF!0�l'��R>����r85�3���/�pQ�@�N��W���J��)����,3��������A�
�c�AǱC'�	�M��)�W_}�/w��sQ���*���X<"+��̢�ЊH���P�P��"�]k�"ڑ`�E������>������L"�w�}ם�un���d�]���*�o��uu5�_������VP�dZOm��%G�|~��䢫�l�Z�u����G�]���f��s�9琯�ݽn�Z�I7T�c�֯_߿� E�0�`�����4�N�����!�� |��8����!P���.
#Ӛ������\iq��W�kGg�sd:g�D%OD_y��K�s��J�(�=���`@UT1-��tKv�@�u�5�ē2�kkk�@,V{S]&ʹ�
�����������nfV��o߾�AzO!#\-R\�Y �fꥋ�&&�AMr�5Kt�0*����װ���l��l��7�+C(���Ckji�+�O�P��vr�����7�Z���?ޏ�'�MM�N��,E�)4O^.G���Vt9)�� lD�1{�lK��h��,#D�J�(&������OyQa����#p��Q��4����M�\�D�YPE�(�v6��e�ꃊ�S	\:$5V�i�fF�ǻ:::D�U	���d]�H�+l�&&R���r��$���U?~��e˖mڴ	t��#C>�L�N	U%\��KN<�D�����!����q3ݲ~5l��V@`�u�Y�vo�i���3�A+2���qzǌ�׮	��6Le%��PH���u|܊"cc�/����0��ƥۖ�p9�y�	W���t�|�_qţ�>����.1[&-v.Mn�+]�E�ʙv��,G~�-�39P����?28�����A��&� r��ښeYœ�\.k�9fٖ�a��+Ȏ��k��Pi�y�b�o����d��^��,���i4ҹ�s�h��y���苶m��+��J� )iS��[�G�٢{-/+'>���N{�"�P�@�./͈�2��p��/�q,��3t�c�d1z���ʤe���4d��ٜ��M癵�wA"bU����'}>3	���@�iL~���r�q8vpn 7~�z#�������E5��AQ�T�	^�x=�IwE6��
bȏnx!��^B������ob�{:wA�o�a5�E�N��ٿ�����/Ers��`\�J	CB.��Af6�4�x"�`tt�@���ni�2�t.�E�V�l��u����S��o��%�t>&l�l
f�m�ٱ�3Ty"�E�������_�z�ao>���}J$�1s&l�O?��J�`�)��}�0QN;��d,�{���<m����a��j/v�a{wm�ܳ�%��8�G.9���ߴӮ(k��L&��E��>g�X&9`��=�V�^->�E�l��-Z�L�u=�+�����￧�rmm��/��bOW\۳�<:)2:�u�V.�fu$J���ܽ�]!H�Q��Eà�͛7G#c~1���Ď
46�I��#~~/Y,P����S��C���խ�g�����޽{���m۶uo���hM�>�9�a{�s���y��&���Վ��`�o�ᬦ�L�������MM4Ʀ�K �r�A8���/U��Ot�o��F_8�<�!��Ң0C���I�B�,��8U?é���Ь��Ŋ��?�U��jH����
EL��d��ĨPM�d���D�\���ԙ>�������o����]{=a2�9a_P9��x�%f��ZgQz�GrPS�,y4]�XԒ��IsU��kj)J��9����sY�C:hbȡ���&�#�SY ���)�x��@A{����ꫯ�f��1]���qk�!0��W�)
>��S�FHX8[Η�s���~�3��b;nʔ)Pt|�<������?�qKgW'ȃf!�ǂ� �����k`h`�$ha�Ҵ �͡a�vP ���)����t2�����k���;n���TVU�C�4���B����᭯_�r%��[o�uJK�9��u�۩�Z����\�{��)mܸI��?�R{9{b�4ug�B�j1���z��B����%��rA�üO@Wc����k�s�}���z{��l)a��<��s֤�`[��@yx,�X�����-�=�������b6��.���S��R�b2�����"�X�G�n���]~�v�����/�ݽ����'u�p�XB8�I~t�U,%0���a�Y��ǒ	��P7�Y*m1S����;E;_ql,� `�bA��e�p�
{Q$2�3��L��1uaS�.%~��I��RT2IT\�@���>�v|l|�y�?pߒ%K�\JX�r�7A���Eۭ|:�
�ʜ߸���r_�fMu��J��*	��N�$Fg��Ws�}{{a��y�2�D����ivt,�T��Ã�5s�B�G�##Co\6[��{��K�넚�a� �#c5Fl�Y��SelV�+�}^*ӓe.�#9��\aO�Ӽ�+�^l2�W|�������Ïqsgϣ:jEI�6B<,sy�.��\Q]S^UM�����W9O6%����,��m[�粒�%(x�Q}T/����C�ڣ}J��h��1�g�,XQ�� 3��ؠB���{��W?���3\"���7�~���l���t*���F���7&�|"�"Zi�!�EG3{�fᬒA2F���a1u(��`N���S��� E!�E�xV�dC��i���F�����p��E���2Y��ޥՂD	��J"FãGs̵�]z�G@�@�Na�c����|�m0���k	/��� N��3fRȔ���윬)�$y�2Kq�X?�Υ��f2)nV7b�����y�4⻠Re��gbz �~/ߠ0(<\,��[��t³2����^|�}�ԋ.�蘣�IC.�]���3�\����o�}����(�(�+���|� ���D,�fW${i.�3��0$��(۰(R
c� ��q�F�q�A##�XC"I0y�����p&P�XyC-����%�����G�1��T(N�Uf���񲘥��$��3���{� M�He�s΁f��������2�~|�.AԹ��@��Z	��eH���֑������J�������	��ܑTr� FL�*qV%����ƣ1���Jd�C��;wwZE��$�!3��	'�R��z�7�`�SJ���ș3����!���e,�u��>T� ��0��t��E�a8�ٹ���l��TZl5��XBN�O��G��#?wy�c��^@v�^O0��g��HL�
�mp�zڄw'�uL�WR��RN�p�Ҷ7Τ�J��t���ޚ����Ej�`����}��/��y�̶�Db4?{	HU�dӿ>��3�C������� ���𝪚:��S1~�f�-��)_ܴ�S
�B4c���H�e�NU�m'��"�\�0K��(�h�p�T��B��`��c`Hj��j�$�S����i�ǀa���uy�tqCu:�Hd<oYN/�k*���{��͟?��?۱c�����:c����C�_�#:�G��yQ��/8]Pj��!%��3�7�Ѐ�$w�'��� �>l���
ye2U)��%%��b�����2�f�(��nY�ϫ++D�u!kj�犳���=;��.ޞ��˺�^_(���N0�	�\A��r6
�K�0��+*y�!�G{��w��T�&���t��o�󞞽���Ht�p9��mM�\Fcs���p4E�=E�8�cJ���l�1:<����J�v��N���y����h�n	X��@�u����	�)��L��D}��$��`���ٳ9�.+K%����Zcc-we�6D��Y��z�ͮ.�~�2u*{#$�1��;o�y�]w��G���g8C*���h���.s�L�m�4��c�v4�bh^5V����a LQSK�Zm�-����+*��+*G��
"(��Z_�L�)*o��q��qy�k/s���I.A�b7���������{�w�q+��{��ͮ���s�����裏^y�� �2��@$�]�u<��.���bt;%�sE�ź��?I%�h��&�'Mp�`_���	���CTup�������`*�B�NR V�%�ѱI�.�'z���j_8�l�r���63fN%Y{�v�-w�܉�(�x��A?M�z��'ِf�����uP洶� z��	��䣖ଶ�+�b�Z��F��W��_�()M�T|
4�8�!K! �ɇ�a�.�εJµ�d��ᐈ'���H �|��߰�ɂD���b�qjj�?���/��<�	�����g�rl�W_x�~������}�p�f͂�rNdD�*�q�n����X�Y'_1�Cƍ��,K���ᢈy}yӂٳw_O����b�>��<�i�o ��M�Lij�����|���w�J�`w�>������_���,\t�ۧN��WΛ7��b&o�R�?��� ���ڍ&ǡ�5��XV$۲<����1������tu�= �����uP/����Pi�*�ͬ�r���`!o���?Ӥ'�;$�#iQ��*R�#��4�W7����C?ڧ̓�w�cY��}�M�\�e
T�������q�E[��@__c}����]0�͖�¢E����=��.��%7�|s*�)%����D6�7���zp���BSxf(�F��d�t�_p:�7o�,��p�β� O���Ք�pQ�]U%M��(�E3^���@������&������ԃg[]U14<&�&u���n����*n���kV�K�=��tX�� ]u����_yZˌ[o����ޯ��*
I��ɤRd����s�ɧX�Y5��&?]z꾮��S8���<�H�#p�L�l౨-ٚS��S@�q=���e�6.�]*nۼéD���gW���S���W���;:N�/0hS�L���p��鳩$NeU�����=,SGU"�U-����t"QQ]=2���{�c��˗�~�i�6���+/���SڛA �!�B�ԩ���'+>����f�k+�Tqf��m�=Y����C�(:�D�u���_����/͝;RZ�<
��:������a�7/��b{{��x�<�������ĥ�9��hі`�lݸaӦM\�k�jFK*r��d�r������m�����?\�f��'�D9Y̑w����;s�L}	�|� %#F��<&)�%ip�pʙgbI�-T?�M'@�˗��g\`�� ��J��j�>�3I���.�[���v��%GM��һgWYY��`'��������I�������;;;:蠎����o���2�r��*�TFw��'㍟|�	�/~��Px��g�jjA�P8Tݦ���W~���@�vt��������g��5���/���d��5�A��q�)�e˖�}�l
�x��>w�ɡjr�e��c7r`p?�%�#(qb�,a�O˔�?����hQ烰q@dB�pv�aG�dgw��/��QY'�����CӦM;��#p�N)�;v�X{��T��)8�յ��)pL�����]Լ�!Xp��n�ԫ�����U���˖-{���J�`Q��r�ہ��7����dxd�*����pE9��a��(��&��>��_�r���`���fb(��
�Ѐ+���u�[���Fd"h�38 ��v8,n_O�믾���R.\�ŵ�FK��`Q�"�Q�F��_q��n߾�'��=���^Mm���Z�~���fL�n�3��)-��,]{�5���_bӦ2�~jTC̨^Ù͚�{n��[n��0`��QV�|.Xp .l\SQ�S[{r82
����d���E�����_Q���L��w�?��; �cQ�9N!�d"���z�)g���yȂ��v��۸y��z���'�&Uk���I}�c�T��h�S�_�	]��B֌54U���e�W����b1b�t"2:<{��3O?�g��{�ʳ��U%>>Q����P-u��O=��s}�_~1_��Yc�(��:22�����t������U+2�dz���㎽���|>����Ï�; �/���C񸋛7o��ο��ٻ��wܖM�W�\��X�e����7bͰm�:��7<�$��T�c����w�ڵ��puUy6���1�ihv������q�暚���=���gp��4�^��?�f�*:T��0�B.�D�d�W_}5�ۡs玃Zs�sQ֜J=��s���lFR�/�w�y�����YH7�US��j��D,N�@9� 9	}Ƿ�{weE�t��� K^shK�xEЕ�(y���y�8ϥp������rÜ�������<y2,M�۔
����h[��H&�PS���wǟ�|�}w͙5gdd���6r�}�ܹ�6eh)I��X?]�f�;_Y��$N]�8�����>��y��ӳ�� Ą�
�΀�p��m$���矿aÆ���p�ʞ��0�8���Ar?���kׯ���x�!P��mm��uۆ���3��4���8묳 ��y�P(6�Ž�B^8<�;�g�m�f1?�:��7�xÖT��
�x0U��x�m�p���$�{z���֬~��;�[o����(>I�ay��4�~�Rj`�F�g�������Y~��Bf^Dp��m������f����?~Ň�}���!bk0( D/?<�x}S#E�8O��~�L���?��S�6P*��JҊ+@^Ӧ��
�{��-���5��Eaْ >�8xε5>�Z��(���=mj�����k/��_��zC�[6W`<UM��b�-��#�{ۏS� �/>��ji���B��  �6�u�;؎�9�rB�[�aC�~ß�Z�����
����?�t>X֜���
"�b��Yg�&:��p���������>:L����a����~�AթN���7�y�i��	'�p饗�'):JؖL~��ʣ�:j����½PPC�	­v/��268}z��!ܨ:���ƣ<���>
�i^�fP�����s�E��@��ZR]r����y��d{�OEAtQ0ʺ����(3
6�ޅՃ27�� �Z������ߟ2�A���+TU��OsO��w߮��>9�c�\!��n��6�jެ�K�.���|����U�1_�̂A]Hے��|�êoo��6�(�x睷-8hlp����L&������GG��0�`�R��@më�y��}�ŗV}���W���ߺy�];��M����~����7o.<"�@+کH�(J�x,�e+̚���.�)w]}��z�6��,�4D���,��m�*�`���c�_~�qY�O<�ͷ�Κf<o��*��8��a.�R��mٲ%S�Zޚ6c�-K;v�%�`����~{�Gn۲�!L/��y���:ܒ$;�cꔑH�E��V=^��KL-k�����9��^����Ν��+��>X�G��8o8�"2Y{�k�,3 ��]�8�e���.Oq�������;w;}��7�,��u5�e�Sfζ l}~W*݃�h��;Je(��-�-P}��"�W9��m"�EQ!@���$�[��^�YM�)x����Zp��X,�����?��Up"�q����:��L;���_~�+<��7^G-��ȗ��'�xb����'R�Xuq�`>o���� Gȸ�	�,L������:U�NEH^���Q�e�[��-�u�Lz�g���Ǝ=f�駟^SY�[EI�k
u9���}��ý���&孌l�̬D0����.2�����z{����(�� ���$��K�~yWY�#*�9W�0L�K.�����l课[	���pb�������u._��Є����9(��4�ׂ�a�v��3 J�0)���?q>+��ڍ���Q\
J��uׁt���z����P �wh����a�Y��3e�SID�H��� 8���$��>�����<<R|����  ��L�-�H�� ��7g��@dvQ�Kv�M&Oæ���^�[�`4�E��N�'$�<�ȃX9Yǀ��	)p��r�ZS�ɡ���hEEpɒ%���œq������3!�9����h���+*Tl1ꜪCaf� �1Bt�����������ڃ�޲�z����h�Aq��<��k�h��9��ˑR���,�'�r�-U,:��	��K�^�(�����-w����倅�Ǎ<��㑡a���S��z�!<�����֭�IU�.*���y3��×;���� H0�ή��ӧ�|Aj�\� �Q�2��V2	���a�?��P躋��b	
_�����MY�2��9�6	t#�����2L��������!��~����)9,ifQ)�[Q�9Sר�8�UWT��Ł�C�w��G�X��f%,*��U=���V�_��g}Π�%AS����:b���[��{�9g&5�D"�`�kk<7D�����JdaW�3�RAV�鬷�͎��*|'v�Dz��-����=;��3>��ө����S��������c���2|�y�J0CYE�{()䳣{�\ud��D2R��9�!;d�]P���A�v�WWm^��=w܏CLgƩT@W	8��fI�74O�n�x6^�m�i8�c�DUC��q�F P��<e�܎���;�W8�-^�+���)v��'y�u�������R�\��7;X�w܆aK[�r}����ސG5T3�,�ѡښ��u�1�q��m�݃�m�S�����N;����ѝΧⱞ�]S��+R�L��db�h���U���A2.M���ܼf�ZT4[MĒч�<g�8�k�|��9��eO}���8e��m�	B���{�+��^U�l�����a��8\�x4���D,_YِMo���|���Ngp{���o!��.ϓ�57:�-���Pq5���GG�������b��\e�ȸ��n��ƺTdx����i�wmߵ����륚đ!��)���ߵk�/�ڹ�����8���a����VՄ���� 7#oɶm`ڶ&@�$�'��L�h�T]E�ƀ�(��	�̘y��!i*5_;ɬ��z� Ovn��ݵN��s�"��f�ٯgsZX����*�1ŕ�઱��t�ܒ��k���(�x��ŋ�I��������0�u�����T�0��!�)���
VQ�JڬU��CTlQ=g��P�H��Q�-��CC�Ph�� ���)���<a沩��V��ҡ�1( ̼~/��c�ǣq�k9=�KePv��wE	��q�F(+(�����Vx��]��;ʈ���j��icc����V�8̩v, !�02�)�����8^��<��FӤO�����rx4�`>y��͟}��k��O�S�4=X�l��ֿ_5w�\�Sj�Z���o�^��g�xi4J9peq��;ʸ\��18�uU�Ys����?e����jNʯ���s��m����8W�c�@5'�a*�Ebb�z���A�f�WT�D������6r�YK-Z�jժt,�t� e��#89��N��;6n܌W�Dǻ8� \�99����6E�~��G�e:Db�;6���fD{�9N�r
�d6�53��,��,'��I�売�R�$mL�*���	�MM@zdL��$�2n��y��1O��D0��fך�A�,%&������l���1�㹹���z�.�JC���J5�~w _(�s�Xti�WKq%7�|��v*9T @�)�m&���gM���_���t:54ا2�*oe]��F�����v���t�����j�[��;�.E��2����\�h �����ã#"J�7��AL�E��.�G���C��ꪏ?�Σ�=��p�e��U�"Q.���g:�c�I'��ja��@�фé{}j4�c]��T*׫<T��
�]u�����n�X)�GuT<���P���J��D�+g��ӦO�t��/>����6oݠ�fKKS6��n_��/���/�!?p����<r}�ҧ���~l@�ۚ��.X0Oͧ_y�I�W'�y�Cmz�wwg�o&!��(\JC[{(T��] z���J��Y1�����ҙk�A@����75���v��=s����Q"�p�B�
�F�Sby,����v{}��_�r'�|�)�P�K:F��T�;��n�EI���~��o��k��A~�A}��w<������类)����U�R��LY8z���;��ϓ7�9B$MP��S�RX�,/�n���j~�Ht������M���� 
2���]*ׯ����8��@�	����2�/�3.�Gti��Ԥ�V!�N��im�~ˉ�Eu��m�@0d�=�5��F��ȡW��3)N��Rɵh�6?��j��G��J�`�\(�5��5Y�j���! ө������S��-u�z?\͊
�z�L}x\յ��ӻ�dI��"�0�`0�@x�J H0�!$������㥓 i��	����c�^e�E�O��s���#%���4ݹ����^���qW�J�!�\��c�U�ɠ��[�Gh��ƫ�ؔ;q�dM
��E�N�IQ��F^02�C�<x�c�ؖ�;o��F�U�+_�dr���dA����/������iPb����ݻ��9��4��%G����V =�3}XTѸ8Iべ��9�Q �[�zugg��Q�:�`�N����%@�E�:�$�}d֯_߹0�jժ��v�#�`���H�
O��Y�/�g�yf"�ۺu�`�9�#�zQ�]���)�2��[��ȁ��oh�c�M-�@�<�`��E���s���i��ѣ��~��_<��ܳ��n������/�}T�X1�B��f2ً/�����D����sZ�c}x��1Fl$	���J����$�x|�7�7W���� �=��aa�:��$qU��iB\�G�&t�䪖<U[9~!J����BuTf����e��L��N�j�H�2��Čd*���`�s��Y��2��@aR}���j�r���|�������4��.Ie�5Y4Kl�-�$�)��/��j�,=�m�J�a�-Ku<�wݵW��=��ϟ7���'��2)�=r��d�6I�8r4��&*
m�e���LMOB�e�x%�H��(�~뭷����%D����z����W��o?}�x����G�5g�j2�T���?��gl����A�\W���!A��4M�����l.���@�z��}�xBP�����쉉����.8���v�ѣ3�'��p�.�JŒQ6̼1���/�p�k�=E�-)���d��M���]nFt.��e��7���D�,ɚ�7糥T���淖�Z��]���}�d@P��^�������"��W�~�p H�C�r)�bT$�	A���GQ�@�Q*��P��t����|�k6�%q ��9�Z�P�t����x۬Y]�ܻ�*��{.$��"�U�O�NZ�p!GG�p,�mll���k�{os,�袵�#pn�c#}�L"�hR�	���$3sOD��I$ &l.M2��-�Z!w1E����*���D%����Oت��rTC!�R�+4ȅ8�&���4����$��A���U[7}~JBҨ#�B�MC��[�])W$E3lǘ�T,rI����b4�܅�)��0W����f�6rq��
n�����{��:�2��������(bh��x�C!��8p`+����o��Yٌ�C�4��x�b�
�\�L�$�d	3��q�v!$���f�`6<��_��WX�x���X���	���/~����d�`/��sL�D�����ܕ�� D+"F��7�۵c�_�6o�|�𲈁*[]G�)k�{^@M�CIC��Ms[�6�.��Ν�q�>��,%?>w�q�$^B������#Oh����Y꬛}	�������iT�G}�����;�8���7�������[�h�'�)�Db�L�u�|�CR���&�a���R�:�l����mڴ	���Z�o�y�Ɩ�æV�!z���eI0|�D#���n|M0�(��Z��½�2_�s�=�]F¿��A�9��3����S����]�Ձ��(���<��GÔ|wd��D�u~��ͷ��s�]�}lǢ�8��U'����0_�����M/6���A� �`������`d�8ҁ{�~�&z�0� �8t_�ԇ<X�AL��*��u���, (*cG�J�i�#f�;G���@z��n��]Y`j���%�{"$b�4��lK�"���x��t}m]cC�-T����_?��<�uѶ�X,16N�,�#�;U���K	2<6Jq�T̂	�h�_Cc������7�_QJ�l��TM�U��@~�ɤ�����9�!�##4��h��5��Al�x&�{ho�	���ښ���u��f57z�O��͚�908�'��Y��fq6 �nvp��x�tv�����aJ�G�ł!yj>W
G�ko��ʧ>���Y�FY�d�(Y@��c�3;;�z0����Vvl��H_�d��4�L���?kƋ/������-���e��j����o����V����q7-,L�P`��#~�aQ7'������t�D
Ţ���Ɠ����Z�V.�-�<6:�w߁�7<3:9��F��ČA�]D�H$��X���lg�t��C/��ƴ!�`!Q.NSKAx�|���;���|T���OeEs�u5E��1�����Ngr�Vx�����N�y��$�$$J�%�_�R,�}�.�F�4�	�N��R,FRQE�
�yJ��lR˕G,���sz�b�f�&ǦYwdl��`D�[(�T/N�@�x�B_ȗ����S$ĤbMT�W;�if��0ASQ����2f�H8Ug�̬�G���چ�b9�y<��{��7�|�����1�U�}K#�_~)�A{{��l��{@0Rq�L��Q��ј助����YH,#��O�E�V?�~�3�ٌ���|*�D)D)��bdU��T���l ��i(dG<������{��Џ~��U��Y�r%��vuuAg3�*O)�*�0`�̓���R���x.�y����O¥�i��n� )���o'1������FD� w'�&�y�m(x���8QD�e>_loo���G��۷C��w-�֐�-���r�����8ls���`Y0�9g�'��3"��	ܾcסC��bwNYy��I��EAi'��D�
�R�+,�� \��<�$�`q��b�̙��<4fxh��E\�:�4!�����,����c�e�`1F���y�x�V��/ȡ
�:/Y���Z�z��CD���*���R��V�$b/L������(+a��&ݠ:]$,lO���,�o)�b�Q��	,�-?KDS�(&�<rȢ�US� F�Q�������������p�%��+�%�E�����[�Զ�6�zX��fZ�4�i|��Ū,�t��3y]�����[�ۚ��I5�톺�񉑱����O|��6,�cf�ֶx᯼����
�K�ۋg�HP�;�p-[��\63�{�<�H��&�b��Ek�X�����Q�pL��0��b��76����Z���z�7��U��~�x�����)�bϝՀ�&j����竫#�24z]6ʴ�X�&79��&�03J<^�>s΂���d�4�.V,�84<���(r��?����w���Jn,8�������ƽ---�᱃�v�À9ءb�
���d,�?��5�wl}��G�.Y�c�Í'Jզ�FG���2�\r][��O�CŊQ��e[���e�*��@�^s��X��c�C۶|�Η�n3��fb�[�X.����4�*�6��z~��	5���oV,��m�v�-UJ�OՅ����6fs%Y!�<6Y&[�dESS�`� ����uҼ���<ϧ+8i�n|�T�4�SG�?��V�&�lnn�D��9�uɮ���ArC��f�X$jmU��
��Bd��u����6Ģ�b�k߸�X��Px�h��ES8�8�3g��D�M��?��X4T.�}x�BCB�VW�FR1{����E+&�)����(f�M�����I$��8�kޞ={p7?��.��E�6���[p���_�fͥ�^�����6��կ~��c���ŀ�����~�"g�5 E-����:�����UW]��k>��*��'��7[q��e˖�w�y�ܞ#�!��=�����D����,��[�E��T�L�����se#_����'f�'�m�����|�I�h �x?`�ITY-��Pd���l$�rcp�Iˆ�Lmv�W�~�P���yI��NAc�~�w���7����a�_ɗ�*�8>�f$�nk��ӭy��akk�qɒ%7nܷoܶ\�Y�|���i$`�2�!$TET�[e�~ n�IpM�S(}�#O7 xK��'%�}��2v�\o���27)� A�ZEr,���X�Ç/?�d�D	��S\�
Fq��,Y�h���G�V�mن�hT�V��K�,������o���/<�O(��z�kp���ְ���%�����d��=������ea��z���~�E"N�9�Is����#!`^7�V�0a�x��x�f!�,��T��J]Y0pK|V��9���a�;ރ�l�o���������ǁ��Tr4��q�@���^w�ş�h``���ņ��A���C�a�u�=���w��'�|h������j䘊p�ۢp%<�?(ҕ:���D6��?x���O]�e����c���ܝ]]�l"�}j���Ơӱx��s��8�v��8�ES}=Q'z�A��4=Q�8�.���H�qF�$���P-5�e�%_��@i���jR�: �"��F#�-3���M�|�P�1:�բ!Y#����:p���'��@4 	 �`4b��������:�
5�J�O����/�v�iu��=��K��)�\�X��t�ssw������]�������i+��w��C�]>m��;���t��ܹs���5�/��b����*+
x�A8�C�W^���>�{~w���G��z�D�U@4�52P�r�H�~����f����a��0�y�}]s��A�Ҭ��د��1k$�IhF�p��0TMv���i�	ɔ���8|%"+YEY����p�g��D�e,��k���.���u��O>����W��u�y'�CD�)�Js��>����n��7�^z��������q�a�오d+bT�'����b�Q�1�52<
	��c�C��i6L�?d�C�UsGx�X��@8x���I'-�?�����>���\~.��][���o�
P�k���,XW_��4�/@��P�%�{\p��SW�NO�z�{l�����= Ϥ��@�b�w�!�r�LM�	|��:fu�%���=
uu�%���\ [�w�.nZ��NM�ee�.n�
 H�^�e��_~�Ёk��Vq��n�mp�Jr�	1lY�������T�t?�Fx<d��.g~8�(Mq���N#b��IVȪ��
�7��:��)�g��?�;	� 0+�\��ĸCuj�+]��x�砘g��cc=���o�-9	j�<��[Zg��s���>�ѕW^���o�-�~����C:���s΁�kmi�f�{�[�z���o�)Y{�ů����ctt�-���]�j�=��l	�F|͢����C�_����R�8r�$���H������<"v�����^���+JU��U��
�wJ�G���Z��i�����'ō�s�=��W���?�O�:xo����΅����~A}��W�/���
Y�s���US�|#�=�'*_ ��pdx�����򗿼��ed�~N*���?=v��駟�c����i�3�кu�֯�<̀�ю�iW�<>^��أ�~��g��E)��xA�����b��C5����埼T��A��ph���g�9k�����7^{������Yq��Y�6�tQ�&�����Je���'�I1
/�X�����C�9�H��J�5�k�a�gS%�����kh���n�v���#�߫���,P4m3�H�}!�t��>t�ɫ��wW�[ꩨ5�1+y��Δq�j�C�y?>�"�J���]�?�9��zm,[D����f��oX�hl�| Q<�(���5�"{���F��Lv�(���h8
̍CC~oY�*"�P�F�2uIu�6���|��g|��u�}6�h `?< $���=�d��/�����hSCG8A�Z�,��R�DS�ڏ_*٪i�G�}������l����MM���կ�<]8<�D����3RT�J�P��3�<a�H����t�W^���-�x�%�U,G��������*M/5>��5��#�b&�PB�S�	Y��7��xC�[V1�ϘѲs��x�)+�f���e>y�5����7�+8H�04��Pxi�-p>����g͙�p�Yk��d,�s�猳O�\�E����x�,ƹ��������>��fsD��͢�K.�dNל�o����%Vo_(ٿ?~�[�ׯO�$����t��r
ح3�?��O>�ԓ�� 9�jn$�q?!s�@��C�AѮ]��G�&��F�޿�5� "��N:�^���K_{���zq�gVG�����7ﺋ)=��^��^x���<��=r���嫸����1ݬ��']]]c�r�$,*�4⌹���R1�?�E.
�[�,BE�F~޼y�B�
jeZ%�O�y!N�L�;b�r] ����X6���C
>���|5��J<r6K�[d1��)t!��N$�*ķ]rĀ]�1��wQ�A�x�WR� �0?Iz�5��z뭖b�K�`�����y��<��?�ְ������Pm��#`��8��[��ŧ�ө�2WX�n,�IU8j�#�,'�׹���,6AQC3M����;�Ed�gf��-�OT�0�_"I.OC[ړy�������j����6��� <V(b5J���_��-�_|q8�|����{��p����$~y�5a���R�2uc���?��#��^lm������O��6Aտ+V@�}��배|"���o���o��P;�í�66Q�����[���?
����:t���EI��!4p]�J�
 �?s-$���[w��U_[G�Z�8x[s�����q N𞩱0H�<n���^���F�x���04�+΄�X߽�n��ȑ����x4a�.ysL���z���Z����F���i����<�)�����?Y��,1DN�75:>I����Aq�]l���G��~||r��`]m���PM2��y��u�L�mјE�Fp-�8�,�4*ԅ�%��
����4�B����P$p\�:�,�/b��[��m��b�.[f�,�N�rf�,���1:049:���'�+���] �ԌM�8�&��=�y��xSZ(�F�Q,">^<^PS���G#�C��N�����/BH�`�͗����+W_��3ئ�?� Y���;?�=␭Zu��'}�m�a�xE8���P���)]�>p0�b��%H��mq�������JW� $1�݃�]SC���8$�b��;B�j����,!���oS��M���&u��B1/R�)YS�y˖�G���_/Y�#�|&KQ4Mɕ
�	d�M�mh�L�7��i����8�ܽ��SV����|��r��
���S!A����o�ZI��+_�\{�Y?��u��������FbQ[������8�3���r�!��۷o4=��8pǏ�NL�[� 9
�F1s���d'F���GG�{�W,Q� �2��|��@����0���ÃCt[*��P_/t�|�?(X\Sw���?�c�
 'U� H�p�R@�d�ۇ��3�6�wZ<�A��1�L\��3�	���`��o��3g�4&l��frU�D�P��v����-����t�����\��p�,��z�Q�͔�VJ(�0�T2E�N��YN�P��-���v'*s.��H�#R�4�����0�������a�����A�iʈ��	"x/�<u�i��#̅�ŉI\v�w�СC��D���=��;JE|'͢��c�D����R�޽��7��>��mY�f�����n۾��죆(2N�iB���d�>�O��KT�hI��+�p��	Û���(%u���~��(ym�\���N?�(��)񩪺7%��txP�я�r�(l@_<��C��,�(x1UNtb()�H�\||*p��'�xf�q�)�`��qU�
�z�ʂYS�p�վ��;�������}u�\A�A���j��� H��>�w�yW�A�n�>`:1փ�{�MW�<1��7���r
@�\���hD8e�ʹ�v�ޕ�f���9�wƣ1��J��:V� �Nd��a93q�y��쓅��X�ffmb0�߿g�՟�������Ur���P�c@��ɄkФ�g��{$6�,[
��I�o6lˑ&�T��S`z� hmj~�t�Vs���s�W���g�+2`�_���V���2�Na��<<�Y�h�Xf"�q��+��4�JQ}�@Q|��ks1�^�c;*Q~+��T}���P�BI�4�����������8?�t!W4O9sU�1#;�2�����W���z��ొY���]��֙݇�/�����x��?6���|�
�H5Դ%~t�7�r}�=��Tm�����T<`�e�x���9R�>�tKKK?,5�]v����[��F�*<r�����f�4�}y������_x�I8�Ӄ˗,�{뭭qŠ!�!��˹�@�z���o��W]�կ|�Lo�)0y�T(M⛋F|��R��l^����׵\��a�C� ~̐���Ԁ51a��h�\�*�IA�YY!���L��>�Хe�ظb�%�7<4�o�U,W�5ǂ�"�f٠�^�c�:K!=v�d�^�&y��p$^檳���qښ'�x�}f3��O�u<	��°�pSe�*U�T*�?8�����/}��ϯ���uO?�\��0|�K>q�L�����2JѰ~�豎��O^v�������a/S_8{����
�y�2<�k/��4J%�\~F���Ev�����n�f��z%Q8�lٲ���D���}�=� )�a�UW]�:�#rXO	&𑯾��֭[�-]@ԋ� �W_s�P4쇖�?v�(ZQP��f�1	�с�B�	�R�G�۷O0X�(�H�H�A3�P����q����#T�
,�ɘ9���!>.�������H.!��B{�f��>3�2�E�,�)������x��-�vu�҄Qj�*W4_���E!�D�|#6H����V��;�!�5)�-L�Q��D�ٳgϻￏ� �LQ���޿��͂���N#Jd,&��j��CS�QWD!n�޳r��x�W_}�g0�� uظ��n@_����N-H�5���6P�̓�>��>� ތ��<6�yй;�1|I��N7�7¦��aP�h�.����y���i����p1�����9��;`y)b92�:o>�&-@.�]5�>>�<yJY&���9����G=e��x,�EX�t)��+�q�!;i\����o��V�ȹ���3�Je���ݏ?���s)�W*�5����b�p�רҵ����O_�z9���3�@�;9��0�?H�ǐ� ����iP�1�#L������R$�Q�a�!�H�خ361M�auc�U�8�c=��o�,�����W�l���ΆN�.�������(E��}�蜊���l�'^H"� <	`<k�
*Ѽ�e��
�R04,�țv.��n$���-��P�j+�BJ��׈��� ��^Q��U�jm�B�?ZU�X�*%�X(2��&&�;G"Џu��=��w�FUM�^���
��lQ�u�P�B������D����U�b�x�}8+Gz��^���:��!�X[�-V/%��d��8
a9n�r���&&_f'H�q�F���L�LY�=[��L����`8�j���L�5A�9r� N�����ݽ��Y��J����wpp�z3f̨�T�� gT'�!nhREi1�DJ�������!A�j�$M�E!��}``�xC���N\q�����\������=5�Ɛ/�MS�*slx,����ġ�z�������jCM���)A!Fb	�ecJn��_H��h��а;w���������W\���/���!� Q�)���9��K89�Љ>���X1�6��*��b9�}a,�kﬓt�.8Mu�B�	S��r��1�F%�I(<֡(����KL��4�h/8�GCB��[L��6���)b��B�������X�������C�k�_�H�(!�s#�*S�
ԑU��Ξ�S77N$5��Ɋͥ���L������P4Ҭ�!�~��G��%�b�0\��_��q~dG�H*��	>.B�)��s�v����g7���=X�����b��h�،��T�TC�u	�4�d&E�5�".d�E���Z�R�]$?��e}��QĈ�{�ㅣ���cMd'b>�>�3r��n���<𹊪-\���J2�����n8H��}'��Y`|po�E�Mը�8"<.1W��s�gzT1z�Уj	ei�3d!�i�xF��t�?V���<�?�b4���ޜGc��"&yp�*f2i�q�G�_Y�
Y6νq�{���������3�`�3Z��0C1�]�����d(@�#�֭{�������k�h$
�n��Zn>6A0qWLsN��b�rSSn���*�d`x<��)E��kz�_�|cNՅs�jj��=�hh�8��#�p2U�}��x�`��dsT�<^$k	� a�4�s����8n}��?c4�۴iS��ð���	G]b��9U����kkj�
:�o�(�¡t�̀�E�!4ϐ&ғ��Ӑ��p='�{e �l�T2[��8v�U��ƿ�F�hw`&����f���:��ȁ���S��淹뒆~���	(��ֶ8�07�J���)��O��(�N��X%� �;���:�R�D*���5�Sʾ��axf�l^$9�agF[��wlkU�����0g5}��m��<�6��N��:<:RL���I��F �L:^O�&��3;f�T�����)�6�X��� �g<Ĺ)
�	3��i�l�+�T���?D�f��ԒM��x
�L8�Dq�;���T1>��W؆1��cdȩ��|��+�S�1�J�����*٬H]}:C��P`8�0e�Jf�t\3ǕHnr�	M���>���YI� ׺D�QO�D@���!��]�v�
��.�o�n�r�i+�:}�w���/�z�#�<:��k��'�{�qZc����{zOţ�ż�TM
�Z̶r�a�
Ͳ-W'��c�c�=צ������,��f�r�Ȏ�vNR�lۺ:&�;�D)����as���~��C��h���j��s�O�o���Dk�n]XS>v���y����N���3�������b�ޗCg���@�AJօk���4P؉PY��r�2T��ڢ���U�c���$��uA6x���,�4��q�),d1�N6YU8�E{I�prQ�(U��3G�'ѹ���&C x�m�0�QAJ���O��܂���Y�ށ!2e�"Gwy��%H���/IC����sV�t��d�<(��|�[nya� .�!+�b���`/�V�P�5����<琎���`cl�%�C�"�-x+�L���h�"(bF
\~Ȏɒ���(CL#�fYޜ�#��(TR�IC�w��D�e wK�+;�t òp�Q�&������s)�0�NSy�σ�9�MaE!���!qo�2����-�D$��y�y�-Z4�X������~����:��?}՚3�X�~�?���@GG�d&�7|��_��ܼy���gw,����Rs�H�t�Yg'ɥ����N�IS��$�Lp;wnߺu������_ ��ȁC����8�|��[n�e)tf��$V�U�����K������w�#4��-�rŰ*v�̙6U�p��_�Rj�c�M6J�hD��4YR��e����P��+�-Z0 '�x�Q��^��{�/�KE���"�R~>j��K$R��6U�.���2��U�_�X�>;!�'ΓG�^V=���&	�-�Qj4�I��-�W(�8�4ݶBm�U${��瓈#�EB*�2ӤH�\*a�Z�u�����&'ǩwQ��wQŖBH�ܿd+)�?$$xM���� �grD�BD�nV��|ב=�T(Lf�h�'&)�fV�FG�받@���(�W�ńՀϨ�++4�Юo��(r��)��h��cGG�ҧ�r
B.6��6<"�7�C�li���H�D��{�y�YR�cJ544���j�w���*�l!��s���BPm3Z�|��o�yWCM]vr+99:�6cF�劃��x&�G��M�yV�h����ͥq���}�͝3��Ph4�a?B�c��y�����0_�����s�mxF����k/������f�g����G��\��{J��Ӗ�~��B��}FC2��445��R�����cz�M�C#�h�#$���
�޽{�|����R�ћ3�8���<U}��m��˸B�:<����XS�2CU�E��۷o?r�hSS����cX�W_}�hO7<���wছ���� ��^�^��8�i1��^�+'�tR<�i`` ��"�Fl��d;�ep�:� �:�JH���XTƙno�uww�,���gaՈ6�X�x)G�4��t2�)�t��{m<W4(�������'O1=(�x,�D���B]����$Q����<8H1�x4ʝ���� ~8J(W&�-�� �g
	�N�&�vM� c��@�u��B�V��ĥi���Q��j�qb���VL_"Sn:a�c˥KԆI�̥T4Nq����'���t�|Ѩ�8�J̷�2���#|O�E4���)�[�7�S�y�"�J��nQ�cJS&�L>ՌZE&������|��?���́#FhH����Y��yL��t����S�D~9ԏ��(r�S�N���=d"i�����7��߆v�⛪���jŊE_|�C���9������9��i��/��)�<TK��2q�4��`
������Q�.
&��î��7�ɚ���zn�l�ʬ�*
�3�0��h��o���nT����l�D�Y�{���c/&0`�;;��ST	�b�da��6�3��O)��EՂ��F������{G�9�s������0��(�r8y!XE7 k�
��?%���@������,>y��}�6%�11����8���*����j���
R��E�E<[�s�Y�r�B��Ʉ�	�N��T�ʯ�9�U���Jh�
���8xl�jkt:d����H��ϑH��V�~���gI�g�b��ؐ� *YWu��OL|p�8CC�P�j��"���zT��R�CA�q�b1?��T.��X8ׂ	+!uEbV?�D+�&05\���|1���&b{y�mSj�FF��_'"�p8��(A�azSD��׶�)�.j� L��7���7^~�w|�<����'��vбWE��S�P��	P�����sHO�C�/��?w��Y�����׶�k�)�D�N��yl�hΊc�`�M����r�� )A�ךL5�q�Y�Pl|,��*:��-g7o~Ǖ�W]u��/%G���S��!X]_ /yɱ<����/��qld�q]���i\������������Ǻ�t��PޮC=�Ӵj!������>��cH��(4DRmc�C����e�d�������\p�J4��X�"7���"c'�P����!b/���ZM��C��k������!m�&�3%9�heA��u�D���]"���g?�����q8�en��Ҫ��J"Sυ�|�"��r�,��n�"�	x�}���pI��T+��]��)�ֵ��#�N(X1X�a����(�#��d*�!�[��-�a��F2��0�|z*�(��@�np��o��u�~���?い�,��h^�H���K��ا�ՖEh���񇵂�����̒�+,+i$�WLP|!"YK:_`mK��*w�V��(S_,�x���mfc(�ޚY�f�(��������n�I�wϞ=(��6D��+�J�Q�X"n�X�t)v�ij�A�H4�)�>*���#q��?#�(0��/~��H�E�
��P٣(�!�
P�?����]����`��裵��)��\:}p�>���_~R�ؼ�"&�QZ.�=1��d$�f�MM��z套����g�^�� a2=�魍O<�ġC����u-�`@���:s��݄�'�ӈEB�v�H�׿�YO��65�Rघ���XQ% X(WR��|����v��IpXd��*�4.�&�cǎ�������闿��w�|}��.�hr$C���-JK����HO�cba���nJłO<�<� ��We�|��eO�J�?!�
&�ZNE�+x�BYV���J�6��6XK��@,�>����m�A�
����u�h"��(Z�J��C@<����Ԁ�8��琣c{FلQ�������pi)l��F'�eXq���Z�8*���Z|=�5`~��Sd��0f��@囹Sql�\��]��<�Ѩ�İ8��֏��B�C����x]Tc���u���R�$��5M��\n��� I��qE�q'9AM
EE�@�	��YG�A`��a�()8��\vά�}������K��������Όc4=��óQ����(g,j����p_g[SGǒ�݇2�Q\�ưU*�/`9^՛��*�L:�c��`*NՈ7n\�d� �{�zaEI���d�����`0L�@U��h�X�M�nݾext�k�r�yCJ�zY�8����C5���K]sF!SQ}X^�?Ss�4�E���������@z�¹Lf���}ժU�Ŵ<��	++�Jы�B�<x���_<���?zOIc�.dE��6+6�jؼ�!�9;�=�*�^��y�g�[���x~t�ʕ�C��Ue.Y���Ԁ��o��_�>ni���T?�l���	�7��s������*���� Wv�-��a�4<XJ�� ��Q��O�AD�-[v��v��!S�,N-��SɄ-[��]�.�A5A���>*�o](�@��/�"�Fm���_�����PD�1�w���;��Qu,,/2�D����7���R�5�~��:w�WeXӰT�&r�S-�)>�F+�+cZ��Oh�rI��	}�����3�N�3(P�>L2�F�#�m�D�f�vu��lx�k�����?������ȩ6%)fˌ'�;f��[�p�ﾋ�N�tiLE�15�8�U��	�.o�����>	$Q�ۦQ9ps"5x|��w�;DC��I���)��#���P�j;L�D&\P1��x���I�+8\rD˲]M�Ce�`$��!�	�[��L�߿7ࣸ\c#�ee�a���K@3�X9��5��������ڲ���w��srH��%K�����@�zU�OǛٸ�::�ة��3ɩ��\!����������מu��X���#�7�֓���!�-�>u|x���y�7���{��S?���C��ϟ�ET�Q[f!�ſUq�N�����R��2*)� ���X�V(�nW�i��?4x�7nٲB1C����e�gV?˴˅"P�o��?�G����1HGE��Lۨ�p �D�*4v�X���*Q�\�|�㹥R�9�Al ʂt�ģ��	��%8`��x5�D��?H�O�lE�Q��ezb�W�7��@Ȫ�t�bs��,�!9�4�ΙD/$1óBCV�Q� �U�R��I.�O��9ў&��_��~��3O	���V��{jI���\�H��tI�m[��>��k��w7*~��+/O&c�zh3/lZ�2��}�Bmm�e��pŲ��r���ϻw���!���V�-�<����+`��������49xd�b�0��Tv2gD��)��nv��RI��H�vv�5�	X<E�Ww�G{��!n��Q�ʳk�w>ͯ��Q-�Ba��
��K�`f(w���#�ׅTP�}kS;�2m�QT@�2l��������np��/���/�|ι���G?�{|��#G�P�z*����#'�6?*⇐tʱ�0 �Zn!�����=���z�q��8e*IY�5�ò�]۶m۽���E"aZDz'��x�iМ?N�V+H]���Z~�pQ��-�U^����9����w���/���(�h�����mۘ�(m����8�HC�mg����ʯ'�9��@��*�+��;�l�f��t�SD�JE.!�# )5�ד�L4���0�%��9�MO�h�Z���0�ł�c��pEKg�X�p�VR����U��W�.�e7υ���D��m�BR��E)��m[[����)NC�J�N)�V�q).������t��'��A��*�V��_��W��5k��� �'��jթs�Ν={nsss)����;�>G.��!y��T]=��Z՚QPe�+�\�2$V���IP�CGG�(� �玄I��ЬO���@�А`�%x̣���
V,�"=�{/����݋�XC�A� gk���G��p@���2��胦m)���F�}���vK�.�����/}�\�:�ɧ�~zr|����������#��ۅ��x��x�B���sU�o� �9���?�b<FO� �o�ٔ�.�@��ʳb4'��X�"@bm})ز��G�d�����U���:'i�@�(nP�O�[�~��H
�#���Cs��� ����/	����s,�Rҩ���f���q����T.Tr�I&c%*������Alli�^!�ZB#A?���$�@��$K9�SOv:��Db�zM�����2�1w=��QA��Q	T�T��R��.P|�3ݾ����tv���@�j�"�P �HR�[�竃��k��d��QsI�r����Ɔx0x,�9p��}��8��,��#Bj���ub* 2M��J(^�������X�����h(W�'�gɪ�/fd���,�Κ�\O "67��#z��~���޾9�g���9��h6Ӻ�+Anxْ`u��[)��T�4�AQ�%�B!	LL�GcT�Z�	��e�g�O!�$�
6F���@�)r��|���NT��D!��$%��V3�-Tz3��T���5zFD���LzDGfq��iUXQq���T� ~4�y��c����������_�~}c}�����v���;8��vR���{�D�T�&/$�F�(:Y��*�{�Il�nH�{���]�-{�o?p�ĉ5)�q]�oTu�s��Z�3�B!v�%PE�#��F��3[dL�_�,���N��3gΥ�^�G����|��_��?�8��?�ԉ\�E�qQJbXy�@9	?�'�:�=���MB�\4�V#C��$���.
(�9d:�5��&:`������8''<���d6Sd��L(x�\D��*u��%���N��qP�#�U_N�s�5H)��$�ID�$��8#	r�a#Ң���ZQKSt
\����SCqS��"Z�������%*𪄹��v���w|t����k@�dQ������"�I�Jq�e�8��'Tp�# ��Cb��r�2安��`�,�Oê����eo�X�}"���,�<B��A�!�P1Ijx�5����T��&���A���.�J ]�(8�3�xFE9HO�
���"�ba�t1_�M�ʮ�ҳϿ�֦g�ـ'"@���4�.�&"չ�i��G�g�ZE��#��J���3[���3Y	�}'Ʃ0%�C���4����*�bO��t@;yq,j��.X�ң�N�Hc_��D�d��}�+:�W0<=�klv=�Z�����x�@����'�F@��U�ȁ�(�����e��P�����E���DT�v|�P*�bX��tpҭi.��\L56�������ށO�W�z�:::�<a�s*SJ��E�&�+�4_����L�t�)��h��g{�\��/��U�ӖK���������[R�x�&��dȖ���(�0D�e�6���1
{��a�)ύX
�F՘�I#�a�jC�L�,W�x,i�M=�(����~��CGw���87�G��BA$���d�ء8QZa��c�Ӝ�H�X{O���� ��YL�=�;��|��6�.Ul�\��q�����ٮY	B>�0%r
E�o{v�T�}R&?��v$��B�DTG��,����ܲv��l�oZJ��ٖ!�*Q�	�2d��P6������X�18V�k��t���ix�Y��W}�S@=���ρ�l����	.6����&�1ΒIc�\+!��tf�͍ϴ�8^(R.4ٍi�We~Ȉ()�i�
�+���� a��5MJ���Rf	�)��7��iH,X �|��w�#�������]w���jWE�
' ��!�<���S*eӭQ�5T#�>X�T��gY����i�̏B���?q�nuժU\ώE|�g���g̠���p�p:�(U	���T(U�`+��H^���_\�v-������HӚ WP�^����4�;n�q��u5T::1�n0�Cb�f�W)��4vΞ���%�=�۳�-xb�Ǯ�'X��Ls�GuC��#�A�L�2�� �^��D�ir���g���c�R���0	5�\Rõ��a�H&�:3��i��v����?��.*��&n�p���W�6��O�3��Ӹ��L#*i<���?�O ��u�YL��( .���b�"5���콛f��$��"y�	�pWJJ�L\��D�Q��>!��TO�۷7�H~�k�e�η�kϮ]5),�y�]�a��W^y姂_4*"��uR�j|)S�H�OĆ*�$0���4�׎� �k��R^�b��m����B��~y��^����n��2~ {*�.EЉ���z+�M����لg��L	Ş=�uxP� 3Sv�D���>��Ï�u�]7~��h�f0_��U�(Eb�d���4%�1��b�
�����Us֒��Roh�0h{n��W_}��?��k_��̙3y-[TK%	go*>$�8-��ϯ�4K��U���M����w�q�7��9���O?��PV'U�U=��;o޼�DC$nj"�_S4LO�(;�!�A/x�X+(W��L��}�4.�1�&9$��F0�&tM����ᡌs5ʑ�PIgr)�����B���)�+�P�bY�Ӆ��I���LŰ8ւ},䲮m:�����������/�:}��DE��b)��ǞM�"k���#Rc��TV���8��FZ#�X,$��c{�o���%�g��Q��29�],dpn����>/�70�W��1�����X.Qs=ݰ
����� ��l.� �Q���͐0���hj���5������|�-�Ͽp-QW��}�����=����ΦM�}�*�
"�ksև����ܺ�U�'���s��O�$ϴF�9/�&���'�t�A<m�'C2�q9r���l'y8��Eq#�b�ō�Tߘ��,�r��JP���L�@4�ȟ�ڞ�+k�}��u���-��|����4"����8P{CK�ln:�ƍ��Mϙ�ɑ.X����^x��o�꣏>b gLL��5}:0�QS1��h�sb\Y�����曮��jH>e|l�����a#�d>UO۲`d ���&����$s��V�B�|�ѡ_D�7V�MVX";�������1�My6U�UDꉷ����AU� h ��U����)��o��I�O��%���e��*�͎��`F��*[�c��&�|i�XE2����IЉ�+\�#�O����(&��P���5��V���ܱ�_~�3���or��z�|^L%!jF�v>�����f�L�<5]�U���%KKص���&���O�\�[._joo��{�'=���|B��3�tw��җ�=����~�,�ғQ�A�p��bU	dfn�+�7��a�$R�,��rwU��:\��!m��������M�Eup����ͧ�@.o��=z������i�����C�����	��D*)b�
�������8v.�\0��ZB��DMSC�� ���9
���/�2���c)I�gr%�P�:��2��R�����1S\�|�]WS[�j��\�P*���_mc��4�� 偡"N(��0��`��u���w������w�u�����Ά��x;�������U%�z����| ����s�B�>�P������g54�S����Ϛ5�P�� E��`���r����ox4G$g0r��U[$��f{����T�Q�cѹERGPY(\|�USߣ�ڋ�)�oz[���H9
 F��T5���r`j�:h��9�/�i��q֚��|�ѱ�(F`���[pZ̊i����p0��Әk��:8�!�Fx��H�������-8���r$T��K�
�����cy�����c/j��p�ˆ��J�jl�-4W�r��hz�,����TӀv��"ӂ�]�P;8ԯ����>�z姮x�g�;／}�|ER�u�w����$�kk�g�|4e]�NŽ]G(���Ԥ(0S������oPɧDUY�Is�T��pq�(�pbp��T�Na�-��� ��
�)5�S4�6T�礐`<�q���À�r��%�-�p�3�sw���S2ŗ�ũ"�%j�x3ϋ�Xq��7����i��?�B��C�����x��1R��+
����^�w����U[_�m�)��|<x��k׮��a�J�R-���&�(�=d�O��@�:�s�;f�[�q�k^|�ſ�����g��
�ɣN�d��+��d2c�)TM"�����@U��[�WŊɉo�pRq�$"I�ߞDuB��CPm�^;��V`��"_���-�c��+/���~#.u��Î�pQ����ǩ|�o��o��ۑ�}��`���oM]n);np�"��).�HS2Y�PXgѡ�-� Z�r�8*[�)���nB0�z��sԝ���a@Ɖ����^�aD���I��06��1�����/��%===3;�ET�-W�_��������_�����©+Wf&'��a��W��#&�y��SϧE���=�d$�����5PnH��ٔ4�(��c!�v�
�F�(��6c�u1=|dd��hh���+�M�֦�Lm-��˄�1	����E����+��/��^VSh�^�EWK4	�)�d[�CoS%�g��(^)$�Д��&��hk��8.#ciB,��K����%����Z-Z�����2��;v�Y�&_2FF�b�D8�\�(UXx��X���ԀH��bD�D�ڠ1#>M�2�x"f�։�>��eE E����O��"] �*��»Ʀ"h `{��!W��^z)�+��_|���>{}{K<U�~���8ǯ9rC��(�s�Ѡ��J)�]b���
���f�8!�u��@�*��=� +�T�D$9�9���>x�{�ڵ��-�R�h����Y_����O=��4B��"����B��Eׂ�[�a2=���N:l����Ҵ���QB4�D��Å^�A���� � Y�0Ns(x�&��@�(ύ'��%��t�(9�s.dp���r9���-���d��F�е@D[S��`7���P���%{z���U��l�\����秊��Q�%uM��Dv���r(8�=⼉��E���SNٽs;��Q,�jꨈb���po�u�7V�X9�3՘"���;�|�ᇛ�}�&�)cX�b��XE���[��-�)�a�]��+9�%�v�%����_��ȑ#<Z��/�Pp���]wxp�/�g0GdKm���}��D�*z�4vi�R%������$��R	����u������Z(IU$w���K3�\b�N�	����ԃ�}��8��y��5~x�t0�8�.rel��;̪N���צ��ږ!��� �#1����((�?����N=�T�`��{���l�/%k�̎���.�����e>oH4J�T�_���|��k�}k�k�I��PES�{&�L���ZY]gR@J�4
rp�	'`�����8ٶ��9)�av�8�C]y���7��u߯�߶m>������}�Gn��V�����ԇ�~Nx��+v�ˢ:�T
�����z�qF�lU�<�8�6�Q�5��͚e�� ʪ��0.*f��	6���A`����}( �'ݲe^�����k���T��0�3�;z�������^r�%4*��gp�Y������4���Ec�H�z�b*��g��A���[�h/49�NCfC86j@�,�n�A�D�E޳{��eK����=�c	ٳ�"�^���3ϼ�����������:c}QFL�I5�ý��{�=��a������ֻ������j�r����tg"�aݺ+/������� 2$9F��+���뮻��wnذ�Z������#I�th�[��v�+�c�4n%�&�'�3������C�T�@�����\GPֱ!Z���p�֜��+�H��f8�	��_�=ǎ���?�ٳ��K?�ӟ����ƛo���܎����+g��v�)�wuͥY�&!4f��d4C8�O��S/�帞e�� ��P0�.~�^,*p/���z�?q����_ח@IVVi�-^��#3#���ʬ�(j��h�P@h�Ed�n��mБQZmmt�Q{Z�[�4G�FD��X,���}߲2+��-�����{#S�3���dEE�x����w��^{�LT|�!� �n$�o�S�>���|���	��js� ��џ��g���߼��~��S�=���6^,R�.K�Q�ר֗�w,3,$T��Br!�����b)�L�ς^����pG5��=&�I�nGb�ֶ����O|�!�������919������d�p�-��˿�	D4�C�Z��S�Х+W.:Y)*�|�Hx��ui/�!�l��7s��3�\��*L�#��`IqmV�s�T���>��kׯ���Nϼ�꫏>�������e(���~�D��~ci�ɽ�N<��3{�z���R������T9صd߾}�\��X�8z�$�)��q�H�f5�v&<)@;!�6�=f?h�����=\����}�닗,�[�r%��R����#����ޖ�,^��K���}����u;�b�j6q�(�J&ɯ������������@�M�[�A�>�[�~��������,⥛�$1����������/~�1�UWggk����7���*�v����_W���=�X�\�6�=O���W�oŧV�>�͇{�+6��eƸ؍tj8ba9�ظ�M7݄���S?y��7��]��u�= �������ᅗ R�H�h�:g;%�)�e������2�DG)Gg7�[P
�W<����8f~ jP`]a�j��
n�e�-��kiIa��������F�N�vaSZ�M�����C�L����Ȝ<#�6h�>��b`vq=.��F�bQ.aW$F'	F����Tke�&M۝����J�b�=*�/�K�NJ(���6�[-r�9.3�D�N���*�G��7~Uh�L񬤰��'�������왓8xO<��g��w~�ƿ�������++�)P��`�!�#B���e�����a%˖u>��s��}�{����
�@*����0`�={�H��i3���)��N��j��U�1
g���z��@����R� ����7`T����c� G~� C[�3����jm��;pR^x� V�äd	�Z����ł2n���
Yǅ�\M*�r�I����֯_��>��#n�q��DK{�ʱ�W֠�����VJ��9�я~g��G���+����w�tO
|�nkk�,�}�]���q䌈�NѨ�||bB|�����O}ꞻo>���$+���I�d�>tvv��}�С#��������^�~6��P�UQ��K�BBP":,I:9{�j��|\�~U8-8��TQ�_�����G7Ú�y�]8���K��'��jH�j�,+b�K+L��h8�X"����ஈ��R�"f���+�(-!�d���l�k�|/�bY�jǕ<yE�V4�q4x�;l2w�B��v����9O�V�@�R���ɐ:�z�x�?x���K$R}}3��R�9Ԛ�(|i*2qY5;�3t�9�����Or"J�6��h��6����/�g���QJ���Q���a�8��k@��0�̆�)�b���"`1\��r�ŗ]����)���U.؈�fs�H�%֒�k:i�O(u���Ξrmϋ/�T��$]��-���jok�	�gɦ���&���s� �4$�Ei�e���HȱT,�Oo�p�;{����<K#!V�޶�(�
EF��PT|�J�=���z��_�%	MUh>���������u�]�&�����h�������~��Ű��Ї �|�s �����ur5����^)W�l�B�|�O�:ETn>s~r��=	�a-d@<��k�.���q�(�._��U����I�BE�D=k��w�y�����6�N&��R�3 
�"EC���w��\���|�[�F�DV��y���\tG;��)�k֬�	J����p���0"���~�Z�Ì���I���x,�C���(��M�@=��HO��X������>�lN�'׻�Î-2�T�rH��f��A�@��K�0���p)\v����Wz��R8��V4h1Ĥ���b�hO��R�<��T;���T�{��\D�E�p��4KL��I|�ߒ�o��\@�A����,\^�\���#G��zrȮ&s�M�9����#@������.�k{g��C�5�;f�!|��B���պd�q�e���Ҍ���4���R��ryժU4�/���v��/�������"���{��S�����:K�.ݼy���N�+�j
4��7���ήb�P)�)*��eg�b��z�����?|b��d;�f���vf^~���ɻ�����i����Gn,�K�g���������ZE&�?CE���\n�@Kwgr���.���ۺ
�F���N�\�cQ"���eQӪ�-OwWw��g�Ɩ/X�`E����~B�Zdɒu���JY�aŤRLxp%$0�&X����M�ә�sbq���;~������V.�) ��2��^�bQ�%yfb"#���)��z�ߟD2
HHҶ��R��H&�6��a�	�x�u%ںz.�|�q
��& ��~Z�S��TQH:�E�O@���	�Ps���ӥq�O~1�i?g��-�sWW��L`�����ޠ��9��YV��������0���t���[����ϖ<w���#6��_��ovP�j� ���.MU��"u���|2��7j����Q|
z?�Hx�&م	�Z�g����FF��KҘ�"Uk����ZҀu�B�w��}������A4C���7��_��I�;� x6����t��s�)�˗/��g�[eg�3
[��ŧh#U�@���R�G��]�g�g�?����G^���:+?K�F�fCw4I
�Bqc�<��1tzH�"v���iJ0	�Fz��3��@�h,v饗~�������,����?��C�}����4KQ�ZqP*����8�JI ���\jQ�D-i!!PTv%/��P�6ՠ�IX��<�)K�l<뮃�a[�իWa3��%c ��e��g^bg���u���&8�'�		�Ki�� 5S�r�z�Ĉ~��KR��d��2�5O�B���㓋�l�a(��2�HY)>�'�֤��F�5y_�']<@B�n��d ����V���ׂ<a��"�y��U4&e���@������̀��P�Ɯq�Y|�_\�z�jH �$\n
-��L7D&�b��j,A��1�y>[�t\
9�k��d%%<CX&�<�������ACH��E���.���-1�K����ND�5J %�-�����N�lK<�T%�x!*�2b1#a��dF�X7�	�ҫ�_��W�\t��5C�p�v\3d��j�"�#���>u�>.�3y��
�Pb��R��7��}�a;/t;��T�U��;:;�X���Q���Q�p�@���̛�(W�*��*�q(�J�	���CK�����*��~�����~��i��}�������bQpC��]�4�t��X���4/��g7�$��D"YM7�]�6�l=������´DI$�E���J�] CK ��_�� Z����4���Ǆ�T�`j$�t�f�`Q�^��9N�?�]��g���v���|�yk- F�j)�N��^��Q:�Zᦅ�f��i�H
�q�ǚsߒ��|����s�2{��&:C.N(�4	�`}"�� Wx��׀�<*QRT@�ZQ�`�,J�V��l�x�J9H3�=�� !�Rw�i��
C�B#����;��>����( �|�����tdמ��q]3�Z�6���L{�4ۄ,C�2�pD�@#�e;�lnV��i�=��@�cf�
G�No#;��ҞJ��;z�Iu��Xш�������'n�T��JH����)��ɩqU�r���N��p��4��5\
�Y�P���X��
 ׮�%"M�ҩ�m��֭[E�⃐�$l��NM0���դ^��陬[��H�ꁂU®�AH5J!�9��[�c�7�1�bQX8ɡ�kdu��Y�&�T� `�!:��g<���0�\��w���xۆ.��'�|g�
��\s>@ʌc�y��q�|��މL|�w�ycC'�֖�n�8@Orsr��j͹��|����H�F�Z���-J�|�D�\�&�:F����퐜:W��8<@L�N���kēB�1y��d��[���ߕ�#��N	�/W�N �\$?D�}�W��
�лx��ŋ�u�ް��NqEb��O�<Uj��܀'��&�?#�;��Fʣ�Ջ��~Sڨ5�T��w�븸�.JrR\���H��;v���'���g���/=���G�ٸi�BנH���l۶���#��7����`Z��S�x=��IE�"w�S��P��C�M��m+�Fl��-����^���!�D\�c��ѶKD��ӱ�� �/�B�*�,Uiwl� Ŋ�9�z��陙s�=�T�nܸ�R*��UKe��i&>��*�JC&f@�g��Fz'�x�2�Jṇ�4�\��	�?�4L�EkkQ9���s� �M����͗qZ�;L� �����䞦t���J�w���H_�Q��MWf�u|tr�����UD�����'n���_�r��@Q�x�-Qqk�x�r���۵��4E��ăf��;���-�-j��I�Z�rM����.���$6&s��#f�K�?p����>Xl=���g�"�_1���VԲ�D�w���ͮ|����Tft,U���/+�pL�*���X���$K��o~�|n�,܆��g����95����D�qG�JS�� 'mb�Sbꙉ������QEW�fg�F�v�Ţ�kQ�P.a���� f�a�P�j)5�!���S䧥�T�\s���F#l���ದ[R���5��ѕiϗ�����#&c�F=6�hi���d<�nmٷoOk[��Ö:�eF:2��Sgj^#�n�����gpyi�������7�w��D�X��U#�h(�����ʗ� �����B8��:�P">N���B�`@:{�u�%xX�xӦM��8��Ҭ퐻ް+фOY��g:�=c)$8�<���f����Zɮ�_��m�����Qغ��|�6��L�KQW���[��'ŦU�0��o�)��UO��>�R?�g�"�e�����ԤO��Vbvjv��e��������)�Ziyh$�i2����S���T�������P�n�aE�צ�ց��*�ºP`��aGa�N�CX����)7=%���'@�/�e{l:815r���U?�e3�ˮ]�֯k��ן{�z
�rɒ%b9��閪�� j��M�\����<y�&��L��Qgv��y���r��/~&�^��H룄p���%j��t����I����R҃۸>l�6ȒB��f��� �w ��K��H��q4�NZP��e����Q��bs\:H���L�|n�2�>E_s%��ݗ���F~E�n�4��̺��M��(c�t!��,���J�9ŰD8��,P���C�q�4g�g6uwP�V9�u�P4K�d�X�@��^\�0;�ʴ�t�K�����yȌF��4*� �و��vlOr?�_pu�|]JsEؤGT"���=+,R��G�*V99�n���?o���3�<s���e5�CM���{?;��}d������Qo�$o��U;a�Y�~��_����n���_xv��́O$��}�}��k>��O�x��+V`OS�����
*:��MPrr(�*'����������LCrJ%�Yp�52�l�W��N;�|��hKc滥B��]�q������H�"Oq�����>4|�ky��ﲫ.�������n�P�����s��/@S��k���4�!"G�x�D[V�iR�C$!I�y�1�x��YJ�{�k�C�PE��Y`���T�V�[� �gϞW^yb���^���_��_��I?Ќ�U�Q�Y4B��\h骚��e�-�cpR�I�����E2��Ƥ�<����j��hMGNk���� �R��pmk�:����v���?0���8q�c����R��+�e˖^{�#��G( V�����4W|�xb��*׬�	.(�
���|�
�3&]�R<��X��"�������:�!���?�{��޾������z%��;<���8��ś/�f*{���Q���n ��;J��'��T�j�\ب��z;��75���k�8�T�S���iB�A}s{D_��F�ON���x$�D9A8��	�Q�@\�a���allt��0�.���nY��Ͽj�I&Za�u,^R:8�i��o��cg[[;�v�����U��"�1���h4��;q�4sgg׉���J~�%��r�˿{�4�OM��ڵ"�L��t�Xqn~��A
�~g[�s��#!��� ���9td�G{:����8���n�TT�t�b�p]j ���Y��d=?�D�G�`���]]�G���;zz:�d��y�;PK�ֹJS�Y��XB�xY��*�b��EBh𠰹c�����Շ��*��CzN�:3_q��^}�բJ%�%Ia�p�\A"M�Ԓ9�j�)"�Д�&Gj)�*~6���яcW�*�ԡC�/	f�?.�+|�c�3��p!����o������o{{����x��o�ۗ^z)�L� �[A�&Ϛ�=&�O�'�(�vX#��}���3J��)l�c,�$��A�DY�l ����NbC�ן���S�v��%���
ez�����?���~��[o���_���� $���0�Fmht@��7R�1���d\_j#%��ԧf��\Q�:�,�K��H*�c��d���8�J=D�=�޽�S�����>�DE�N]��'&fZ;;H�Z}!��Wd���y~CL�|[�'d-\8�%%
�h����8gq���z�a�x�����X4��;6_��f��R�$�����T,s��V|��ჿ���! �@!��R�4���FM���C��y��(��,]���8���s�i/���U����3t�T4�Odj�PW���y��;��x_G�y�Ν��Cw���C'N��G?�}���[o���g:�%5'4m��t��y+*7�i<�Τ1?|Vq�=���?���F��I��H��4����ߛ��!F�����o}�8Y�T�RK$�\JK%u��R�s�5���w]k�*�J_4B�sJ.��/1'*�}kY@�Z��R�rCPnx���'�����k�$���<��y�'�ez��a�2�~�a�ՒS�ٽ{߁�;a*��A�fc�X<Ia8��J9_�bG�x"Z,��5h�e�!�C��Չ�<��b@ۓ3��J�Z)��y������,O`������o���D���g�iR����.�����O��oX�r�¾w�^^��x�".Uө�W�E�=���9�/Nce��\�>S�Ն��RSA�Ac�������s( S"s"M���:G�L˯�*��[M=���C;eW�xB��G�^Gg��+���tZ��BaͰ��ݔ*�U3�
5�ˀ�@u���h����(L�S�K�v�ٓHF�F����}�5t����xq4�Z���-����[s��L[�k,���"�Ru���6��{cc�^x�ͭ�vfG[�����!$��сI�5��-C]�x��%�����3�>��+�}���F2RAs� 
���/_6���}O�nӦ|�P�۶m���-ZD��y䝴ۈ��������w��&�-s�B8�g�b6���}j�:K�o��W#�	d�x&�'g��f�dǬ��Ee���غ8~Ŏ�3������(*'߰%�׺k��֘泌u�u׭[}��c�a!�6W_�� 9��wދ/���XO�XI���V���'>��x�U�g��L�Bա%�b��A%�.$��B�"���*�$u�)�z'�1��	�(��=��Ln�Y�\f"U^~�eέ�8p�[n������?�_۶C�J��p|��pdtt����m�'�7Pp;�$S�Q�:{��SRY���#�{����S��}f�OD�p@g�k���t�b5��h�)w]vS���(UzE,!\���-Vl)Q��@��e.*�5�) �W�ٳݚ�0!�?�� G5�"�W\N� ކ�do�\���ƙ�N2��ݛ�?���#����F��=oc����Vl��ŸIhmZ(����Z[���_{ٮW��
,$��׀[(]{��Ν;���U=���!��ݮ���������O:�/;��a<yfA�׾��E-�]����o���	�.��B����R��;���>�P���ph��lou�0 w�+Pb�Z���r�֨-��yg�Nh^]i��X�"]ˤժ��4P}��6P���	U��]�i�3�6	��琅	��Jc|��<P�+W�������É�3�H1��]E)ը�%Kt-�����+.�ѹ˗���y�(�躵+����N��L������R+;%��V4d�׀B����8�Q,�].j�p8�����ao�d:�T*\@Nߞ����r��g�(/��q�^��
�嗿���?�ݓ9����%�]-w���?�E��R0:a�������UM�dg�P�!8�ф�)�BI@ ��@:��]r0G&)[,�P���sEA�0)���'�*!��*�+P� nm8B'N��]�:�����TƃC��ކ��VG�q�C�}W�7	�����!����_B�V�f9���]wݵu����?�Ꮢ���י�p��~��m&�+��R�ACC�ȧO�����zk���K�P�A�2���Ⱦ}�~��ݻw�n_��o�N���㏡p��hmzQ&����׮]{�9�P^�JM�CCCP�����JR�'Z���o�3I[�Й������f�����g޴i��7�!d�B,-����	��yIa3$r&	=,
����ܻe˖��V��(��H���X�/#�2@�+���N�Z�&���>��CR+�!�
�5,�ӡ��1���f~x��j�[p$Ն��#�r6+���@��!|u�L��L4@"޻�$��]�ٿ};����^��!���W�z����j1����Z��J8��i<J�w@�S��$�j���7\^��x���������L��@��7��������7��|�+?p9|�o=� �^�MK��@��gN\r�%Eׇ���x�aC2���d� �
VQ�dU��@D_��|M���r�FOԱDG�=a��q�9K��|qbb6OQb��.��U"w�U	��@aai4��O*�*.�Te�M�'���CF���5H����ǚ|����{��k�Q`�/����w�}/���l��l��V*g�|��d2�t��X@������*, ���D���%�q׮[�}���O���^�~�E�dQ���ڎ��%<C!�VܮP'�&^���f�S]��<� �*T��e�ʜ-����K�z
U*�HCp�Z�l��"
!\��'�]�x]��<�g�E��cc�3�VkL8�B�W�f�@<\�V��6�u�pv�<�
�
�`	�����-*��f�q�4�~꜍V|�â��~M�p��'�	�D�X(��f���9�2r�HG������J���[4�vbb�η>�����|��������?�q��K.�h��#�G�!�������r�B��琒R�Ճ��+�>	�:�teZ9`���Vk��b�82�Y15P�5	�D%�q�e�  W����Q����ɨn(�������1+l�Z��T]�|��}4IF3<׫��O�+�F�bwu����?K3��ͱ��+�x�H�;G�1dJG���[.H����(��{����	.���֌���H<�?�n�jS���-��9wE��R-S &7C�?cg�����k�20y�v�p7�<	��SHC#�Ru~�\u��=�v�y��|��T�[�NV5Bō�.(XX
��E�ah�$�A�������cG��-TO�J�����C<�-�<y�k~�>|�:`A��ko�_0>5	�ҳ�OH 3\�7�"�â!M�>)�PX�2~&-��S*���T��T�)�mϷ�K�K�c.�x)N�h>Q�T��$�-�x�,�w�J�:-i2��XX�T�¦Vg��U��'��$��CG���n��L�e�q��점T�8Q����T�ȭ�<t*O,�f��Q�G�Y�����E�������h��k4z{{o����>�O����#�K<��tK:�s>$0H	�Lg�?=K�!����ZIT8iF���w��"T�e/4�09=C�5�_M?��͓!h��g��֬�Ҍ�����n�	��j�x���;v�8g��2Aβ_��J%�jj�`:Y��")A�{+:�WJy��U�e�aRr4��Ѣ�fu���I��#�6ˌ{m�,v�I�(*�!3E���5#�E\u�#��\���$ό��{����L���0]���I���q^x!�!���ge�MU5z+�R�a����x��F;8=Y�W���n\`��XC�TŌ*�r�W��w���;v �f��aX�sS����sa �;�o6��p��b��cs���k�j29OnV ��Ҝ;H��gZt����(pl(�C�
���qh�KC���W�6�x�(!��E��M	���\�.�^%���R�%%�p6�������j���u�nФ�Ϻ�X�I��E�����I��N2���˘��ɳؽm[�^}�Um��Ͽ��zԍDbkfj2�\���ղ��\��kԪx�?��**��Y6������,�"]k2��]��E�J���L�M�yf p��6�@C�ӲC�z����g��D�X��:���KK$W�P�j�B��PێKi�!,���|�s���@��(�fg- v<;z�XDQ{�z�a�=�����o�u�ݟt=i�c�|mxt��$�<�M�R�=�<zI;�����j4�ؼ~{(�YP1<�WSZ. iY*ʻv�--�G�N7�4��zؘ������)=hF�[��?5`<or"B�2%�8��$����͒�@�:~B� 䄀��:"DͿ��o������T"�� k��&W�������[�.]�ď�_�jUK2���l%�TC�~rwL���>� P/L�P�A4�-O�jI� ��J��~�R�Ǌ�#5�y.���e֩��1Y�<����vn\u(=�!⨫�w�IM����F��*�f}��&%ק���<��{�ijJ!��h��"4+E��x�n�C2�(w|SU4W�F�禅���F�j{a� �^�O|ꊵkaI$�%�#����ڲe�:��[pd��Ǥ�t�C��.��:��ʸ̺C,l�0qZOM�ߘ�y�?��ԝ"�K�4������P]��rҟ��`��~����n��F�##�z�jh��,�0+��)W�$Ap�S�N�Ҷ�t�9�0��T�m
�#]��(O��8,l�����H(��+� �)�2�k~w`���wR��z��y	j�*��DL�ݡ�mcAO?I�J��dV�SV�Z���r��؝�E��J����M�OP�]��a��,d�`u9N`�t�Z"Q8A�]��Z�C8�睷.De0�aB��� ����U��?��G����P�E4��їP��+���k����X-��\W����C8��(aa�[����K��L�H+g]g�^�&�)ihf���x��Ҩ*��,g����I1��xG�8�ק��TK�+<�T�-���W��e2���|���aa���������/6�G�z@K�|î�-�����FFF^������ X��z�="�R�zgk+�ܙn+_�����^*���xn�xjjl2�Rɛ��TO)���T�D,
�P=[�Qe�|{X��x�f������t2���f h�?��>�Lvff��Z�hI;@~ݞ��G���f�A|���s��%Pf�Bz������,��-��=�'8���)c��[�S^T3�OS����CVv&�ĀΕ����X4Fj��D�c9�RTH;+b�Je_���x�A��ih	��V`�Ca㐌�!��т`�u�3`��%kfq�V᰸R�!B�ex(M"�%���2hX�����,��lQ�T`"����zϖ�O�v��?>I����D�ʉx�q����;!��\���`]��(�������V������}�xc���Z䢊����/��6#8���7�$�����>�&��~�N��}sl�17Hx^[�kqw����ph�5�t{{���8t�=�#��5�^@���֭[w�=�;1Jo�����E�|*��¤�Z�N�uő���\���^���V�h�|���M����qː�c'�CU,Y�k�K���B9�rٺ���I"F� H��Çi��Ę��<[��P(cɬ�UiF����޽e<��-i��t^=mn�JF�"b ���������m�Ҵ��(4�2�i752�J ���a�v��E$g �"�S�"��v������4.�O�ƛ�K��Hj����u!G�� ��5I4����}��6��y8���qʡG��
KI�f����h���D
1#�����pE�7��7�usU2n��"���x��乹�tn�|�EN c�4-6��OT��Y�JrI%[|�*o3-�j5���7������'Xm�~*2&�=S�&9�Um�O��+Z�V���~zh(��/^!w���h*��G��g�����C���Zn�!����cP��ӓؒ��	{P���6�:;*$�ڠ�D���������bP0&#����4�['��a�@S��+[���$�TY*�����I�[������Ĵ�UV8��g�g�}6v�|!E/W+�-T�o�
E��U���x�R�*�0�y��l��fG��B3L�7�@i�<d��������q�:��TC�}�Ƀ�7p�V�����v���,U?�"�����H�I����uy��H 
]e7�>�G���]��C�v�N^����٢�3��d(�杄��K�/������p�pȱ�!��G旿�� H\���ڇ    IEND�B`�PK
      RZ蓎�ɣ  ɣ  /   images/b240e25a-70ca-477b-8a45-be7a3295a83b.png�PNG

   IHDR   d   �   ���t   	pHYs  �  ��+  �{IDATx�<�|\�>|{�>�Q�r�\���6`��I$��M6�$�l�.lvH �M�PCӱ�n�^dY�d�.�������w���	i4s��=�9�s�y�s�2�O>����;J����4Ϸ������*�(�L�u��5ӱ�2̚�ܾ��w��&ϸ�mI2_S]�x�s-ۑE��h�4�fZ��q�rh��8�����4E��l�r]����(ål�bi�u�e5C����f]�ь�a�j��W�M�w]��X�r,�r�I4�����\�uY�%�R�#���i,/4-l*��t�Hr�#в$�65M�]����<~V\�Mq��d���7� �
�˥~��?qln[��cc�%���������%C��⯨��w�7
x��yb_υC�R���Ex���w�	c��\ڤi�r)Ӱp��1.���(��hƱ�X�1L�ʫ�rm�`����\���8�/���p�2�R�8�:�ڛ��$�˚6l���0|4/��Z�eO��q,M�:�ӒD��x۶�ҕ��e�%%��\��@6���`�k��gS���r&����@ �z�R��<|���z��G�������}���JY`�����>;|���++�W_}�uxמ�?��[w����5����P�NdK?����8c#�����Q�ʶɲ�?��u�ւa`/˶��]�k�X�����ض�2��8����1�´׶����Uk9icwh�P(拪�H�	�`�b���-���jÔxƲ��M�����!��Q��H�����_��_��+/��BMU����+/�Ɖ�mw�q�M7R��Ne��_����.Z�|Ū��f�(��j2�:q�L:�z��W=~���:;�
"?1>��{�~���f�ym�.�0�_�Z(�(����]K��d�zNa�4ϲp����<���"��;lx�o&������s`<�?� h�0�CS�C!��PvٚpS(_����S�"�ڸ��ٮ[��,-\6F.K�#���qM��n�0��/}��uw�r�����W;����/���l��;n��R6�
�ʊ��ꡑ!ڡ�lݲ~�e>����F����ς~|u��6mI����;JZ)=;�y�L��E��wg����	lᦺ�vH�x�q�<yth8���@E�5)ǵ-&kS.b���<졖
�EAmX
�`���1����l`��f%^�P���l��o��G��N3���]q�������Hm]Ϳ����N�">��i\A���]ղ���~��b����^�@���[�bY�W}xr,�M��rC��'�����vm2��*�{���hwd����kϞ����w�X��F�Hf�@fQ��(}�ʐ.�:���G�m]����<�V�ExA
�<�O/Y����;��ϩm
+��8\��f�yd��jl��UF1�CsZ�`��)l�$I����z�~dt����QUU�s}�}�|�7�X��������Qhm�x%vh���Cǯ�rMe�RS.�E�`k�E�����XG׆(w��[.%��d㣃�/k;r��2���J���^	�:��QU�����_���������6�N?u.�Ey�oO��vu; ���EQ����d��ũ�˺MmsB�*M�����Q��(�.U(k��b㍍ͱ��a��id����9� 1E-�"���	^�����Ԅ��F���îeUWU��ffg\]��au�B�C\�uqc�=�Pw-r��^�*o�������!���~��#��"S��]��������f���s��}�ݷ�k���Z�e���3��驩�߼e�3g�>q�ԍ77p�|~dd��ݝɦ����8������U���� 2��3g�cct��+Y���Ю��w_�+|����^I��1�Ҷn�8�$Z�����^�.45�G�����������"I&G*"Q�R�P���V�h�><<�,�{�|~�B5>3�9�Vd	��?�����o��۵���BJM�N�2��Ԑ�nmj�Xm��o��_|���^��ܹ5+�-|������Wl����D�̹����{��Xv�Cs�̙��z�oϜ^t�X���|ǅBA�E���
䯥+VI��Kg''&o��@(T�gw�x+$�w����qv���^��U,L�����������z,AY]-i��������9��۸q��ب��.�O"�hm��455��R�i��}�`����p���g�m�m�Ń�V��,5=�u��nᐿ����o2�]�����B>��S�ǲ�c+C!=�7f�ږ���v����~�h���n���m�ﵗ}퍷kkjgc�s�ڐ��������80���ؿ;������yE�p,����D�p���O�l[��%I��;���:��<�x��K}���p8�����&ŐFP��#��-d�Ҹ����2J��ёAAs����j�3��gO��t��t]SS0س�������f�
����Ö�� �x6��R�d:^��>�6�lr0>3�a��x<fk*ݓˌ)r�����4�QyG��[���n|����;B���=w���A�_}�U������E0���5ST<�(WWF�SS�ip<��1�*���}��'5k��L�8���4�2@����ʪjIP`P@,�J%5M�,d]���KE`�HWgW��_�pq&�F.��Z�xA�$�P�)�
D��"��]�ܓ��/{|�e��|��@24K��a�|b*	׶ջn"[�
V�fҳR�<˫���bU�8{vG�~� |V�Y!�K���F���F��B	�W��J�2K�J���W���¹�>^�M�>��? 
��?�������?���΁��'��=ߖ��UJ�)K�`$���|��,����ŝt|�����]�!�JPH�!������Ų!�l>�eN񷯺"�N��Ap�������A�����rL��S�z=~��,f�:(��2"��p��*S7�;��TSe�|�E"�ڌ#�^I���eI�}h �,}���N��~�_UWo���y�Z^{�����.]�~�WΟ�8N��[O=�l���-�믻�*Bޡ��/Y��g�k�+�ɸG�3�Ԇ��O����,>i��yy+q�7��؏�HD�q��xQ�����#dV	�(���1���u���@�ã�d���}@����t�\TI����$��[W����1�ϥ���Q��i�)�O��&����Mkj"�`^�`r�B-��[+��"�p��h�iB�l�몺���������t\EnG��u͛����l�j���6\����at|�y��?�ﾱ�Q��B�15UՆ�&��|���M�M�ʊ�X���Cy�qc�<Td^��������K�ǎ4"�D%>=<�c��vu&��)�N�3�\NQd�
��mb'
w�@W���k�&�/�e�D�h�M���5�R�������h*��h'��j1a&�N� p@�LFSU�q�����D�U�)�567���`vj���VM�L�����-wm�X�<���T�a�o옜+��K��b���-%s��ZϺ�k4|8^71>�x���Ý��`�����l�缗oڸnͪ����=����}�,K���B��Mi�����6f�S�f2����qLM�-�E �c�EApl�Tk�=�	�� o*�7�P|� `㐪�N��%L���D[�������Y�aU�reB��?>�i�FN�_}�7�N�?p���V]�z�쭥$��
���+BZJp�L�#�T#�~��:
����~��;�W�FO�:)����s��ë�֦�Io4�!i|��C�?�v��윹ǎ���@
�;�r*�ٷg��� �TE&�=y�xz&�y|��I�K�������TI��<D�.�3"\��I-���K���&:��$	
bH��X�0۶L���8��r,�Ah"�m0�C����MȒ�gϧ��]ə��/��4�����Z�Nd���i��={����K}����^�v<�^P���B��Dn��M��<��׿��"h��=��S����[��ej�$��__L�K<ϼ��KaP	�Ƈ�C@B�u��1M+�"�L�4�g���*"�U�^�q���̤I[�F+��ejv���nrr������u��Hc}���8���*d���0j�+�b1F��a�`��b�3���#�S���lni��=LMO�J�p0����.y|�ήK�ݩT|�����OȒ�����s����x���!2���+�`�PR�edS�%��w\�V�M�����'���ڃ�OScM(������]�x�ྉ��HKC��������k����hԁ�{ʘ����@\��cO>�d,6^̏4E���W;.���p70�k$I��gff**�3�i$�x<N*S���	�Y�-d��D(ʄ �TW"A8~�bS���dޤ��K3�D��Ւ?�������(��.�t8�e�\�����ϙS�P��{����&␳9�t��ǿ�X�޴�Kw�o<��_�9��gMۓ�t���>E�8u�����8��y��� 10��p�'͘�ٲaC�eQ ��r�ѵ�#�#* Y�E{;�y�IdC�"KWͭMݽ}˖��������F%�G!w�����0R��TbRtffV-�c
��ձ�l8��2��%K��⠝M�bq����ܬ�E�T�H(��2�̊�
�a��"��DHN@� %@�im����^z��|{���];y�𹹭�H;��e�� ��%�$�: ��܈#e#*\U8 �ʤ�>?���鰡	?ph�&ѣ��lIK�[��	����9`�@���!��FF�k����d<�:/O��dr)0%� \X���$D3E�u]Dn�%`��'������&��Z�ZAnl�S�iz�������Y��d
��fh.�	{1���]�)|�QYN�ɒ'��.]�xBъ��=�++�)݆�=|�X"�G�g�Y�I
h�k��@[% ��z�M��D�����<��33q�f���W�X�d��}��?zd��u�����!k���/�Ny���ڀe�]�xI,������D:�oh�C@����dz,�pz{`�	���|mmu���,������E�����rkks<��'���\��/��3�>�4u�_0�A�=�b��'�S6҉�dij��꘲b�0��><2>�{tz�ޣ��d�Y]3V,_�hт�?x���������~��ś7o��];��t�Q��˩��i�֛n�]�����֛�ɼH6�����ܳO���R� H�E*?�D��[o�1�~l����E�Ł،˰��,�l!��==��OMí�or���02�|��%���� ����FЬ-\��<�q�2쉩	M-Ŧ'E^�Ǧ�㘢V QN٥8@�I�*��	ߢ��y4)�;F��>�h
6VӍ+6.�����w^�4$kDɴJw�u������Ã�����m�d���@֮]��}?� ��V�����1�t���
 JK���}�u��}�!w��<�{��9�����8�f6��ֵ�E�$XPI`�&�e�$}�TJq�DS�6���z G��7ClҤ���A��T�M��8��؉� ���,Y��9HQ�����j�: �b\�!�}�hH�nD�m�M� �^q���?�����S�D ��o�����3��6�׃�o�v��¡�()OŵWo*�90G6��(���M665���c�G�{�?��ՋU]SM��a�S��M��$�6ΙJ���H |-s��K��kE�-*J���159n��
�8�Y�����9���x�W� QhQ�'�ܔC���'�	R�'���3��3L�0 u /����������#���bA�i
�ʛl�p���U�4�c��>_�����ܳϙ�0ۭ���'��l�������l���|�����oݺ9��=w����)�H��O=���Ԍ�(�(0@�v��t����'];�y�)�:H��k�+�&�FZD��]�V��d1�N��Ӥ��i��k�F��'I�!��7Zv��><>���pX��\~�(�a�B��Jh?M�".�Z���mX&R��_�K��N����C�_[c�{�-y�B\\�m�����W��N��|��_z���uٚ5�+�5�oߩ�n����?��Gښ�K��� NX��?����V�ݳ	�X�:�n��ˊ�]�VY�$9Z���W�*�u�5u]g��\"���K�,����cj���u"�1���.k ]�v�@E�A 8X3x+~eX�`��$]�k4�+M��4"�4I�6"a��<迁�u9A�MA�Y0�Eږ��3�U���cG;@�DE����?;44���SS[��~��S�T��kh��w���.]u�IbAe����0�X��?.�hb����ʢ�,��!�п��/-7�������h�n;�`89����i������{�mIbw�"��|�'�P7��!F��i]#�Y�,�����X�0�U&��6XI�E�K�A �t��!�D0�&���p2�u���_����q��>}�TXw���r&�&d�f�ώ�8q��#-H���:���,���Z�@��G��C3$E������G>�e�s�8�L����q
 �b���0�R�̟�H���SIF�"ɰ�K ��bbKbG����g�d88�i�L��Ex%�%	8,Ŷ��vI��tp����@7�AJM �N��-����"�5�p�7om��؉���>"u�$��M��t<���e-����)�D���D\Lװu�m���x���I{eqr��+t#U���9��oB�S}2�@�� 9QNCC�6��E^��# &��%E�S!�Ѥ{M�E�{��L�0g��!{�H��8�V-��k��MD�%Ē,�uEg�Bp� ��L�=����m����������f2$�]�P(z�x�X̱�Oöd��<H���|q�5׭^�r��gfjzl|zE �LD��[�ww���<5����G�yn��p:9��Ԃ6�*OMOO5�[���<2<bO�x<V[Ss���5�A��X|����!ϐY�O�t�\X������a"c�_�2���w0�Y+�h�"3	j��D/��/�bʆ�4������ �o����:B���-���o?y�$9�=�]UmXҶ~�ڀ�߽���=��ٮi��u����r�t$�{��Wt�o��=���.���������Ȼ�n!F��? ϼ��-mr��b���ƽ����Kk֮�?o�ŋ�|���u훮ٖJ'��:���3Ij��#8�QĔ{� c��&>b�!��ʰP��̒e��#�Jp��e����:e��)�@F�a`f,��x��do�*�,i��ŗ�^}J>�O&�pė_~1�����@�6l�a��5H�kW^v�M[����r��`��RI�D"�q�TVV�r��ÿ���}���|����g�
�T�}����޳�[�<�}� bE�$H7�ٴ����(1��80g��,!t6����k
/�I)�#]�X�bE|r� ��\*�`�0|~��2I��A�K�"��&0+��d����|yH��-O���$A�[��D�5�jsK˺�_��˟�����g�*���������pkk۱#�V�^~�����-��h��}G&_�D�/�f�����qr|J���ʺi�R��n��-�]gϝ<y̱MN����\!�%CE�.��e�s�I�g��Q������].�1"���|(F�>$����JD��11cÝ`�@�>�P(�2z�3(2f���-W��4a�P$O8������x	�h�*�@��+�ZVg*�+��jj'qI:2�Ҏ7�Υ�`
�2Z=444>viρ]�o�RY��p�,�߷w媕�]{m6����|��wp�إ���;����G�����k%�e��9R�Y!	��!g1e�	��Y8� �A��\3i��\� �(ʒZ �B$���n��$������I���4�@�` �a���"9�;l��v����WSɴ����)l�& IWf�ϼV��	��Uc͚u�.ߐ��v����}�|y��Ů��*��xkǮ�n upJ������O]�=�9J�̿����TMu�L<�D�䛾xcT�C�19�	��b�%�w�N���L�C5��6��bXU�J��'=AB�#����ۙ�a��݅��@�K�@T��L��p�X�%�8]f	�N4�]N�xڄ`�
�a���,2�o�頬�Ƨ��3�o~�Dנ"�q�/��ԩ��"���B��;w"�o��f�����v|zɊ��un I�9�rQFD�!�E�7��ih�	"~y��eꋷޡj�9�|�b���]EM�ˎVV{��@\����� �!}�R�	E4���B����,�X6��+US�~_�X@��G \����:0��Ԫ���4�),ʕųC$r��Bt8M�?QQd4�g���L�+��C~�2>R���fo߶�����{tzdz&�������O
��$�w ��w߾#4o��&+Vt���]��a#�r�E�DPC��%��0LI����N�|��`M���R^E<�R��s�T"���?55��ad�Yo �R5,0��{92��y�G�-RDV#�<:�&Rq���� �9W�K�
I&1{�Fp�%�\BP�k::��ES��R4�0\�um�'b.�A`ݍ� 
����M�zղ���_���rK9��e ���IH�cE�K�ؒ�a�$�!dC�hF	�A�aI%�#��<Kf�����y�*L3u�ӗ�WyDVQ< o6�.�p%�þ�@4t<�k˂�HJIS<��Spr��(�"Aoi�����!\��\�-�D��lZ�L����3���l��b�!�#���������eyV��7]ӰU-ze2�����4��	�2�#�Ji���x|�
P�e�6@��+�L�G�EV�I�K�/X�i��Z>76>���7;3+K^�+N�Έ�~ �q�χ�޹k��:e��cV�2!$�d,VȧD�C��ufgc��!����/u5�֔4����7����W�����:�O�j���pO	�$���Y�vB��ll�V�eA��/BNIo�hI\�H'2HA�R��$:�2���(Wg$�.+R��vf�������8`���H�&�.NCs��Ƞ��,����]�`���W�Nq炙T5�QxҾoii��w��N&�)����~��������Qx�����ox����S�ݺ�Hq���Y��X�\�X���<��43>1�'E Mb�g������m���*DQ�D���rM²�Vα���p���! �
 J�ȋ����R��|6Q�ςZ'��2��� "�H�&i��FX7o���7��%S�b��'~6<`F"����Zcc�>��
O>�'��^u��?��o���kj��m��G��/
� Z�h�����:��o��ᙙ�T6��޾V��W��w@@yz��&S�c�έ\2�ȹP~���0�r�� �64i/�y#%���h؃ 44�� �BL�{5	/�-���Ѡˉ��?y�j	�5t(���L�[�)P-���6�2�r�}<�<H��j�(����H���u�e��{����_�����Ͽ��ܺP���O�S/�����w]8;>�hi���������%������~�R!��­��G����[�y�/S�c�$�p�U�Z��OD�#��j�D�Z�@�g�'e
Hf��I��Ҵr�Y e���2�ᭈ�0y�W�-N��\9��=C��˗������X*��|o<�hmj;�c��ޡޥ˗������M��/���Y��}��#zDQm#s����k[��yEo����>��B����^T���
	����TO�`pU�"�9��9|��u�浶EB��������e�^����������}?�d��-��	���j�7�L�5 �5�u�9$xIf�H��uY���#*��B�)�2��ȲH���ƒ�$B��d$I"<�h=���F���Ed(��r�`�����"�%��k�/^�h��灏�׵V��x�����9qdt~.�4)�9"L�}�]����q���~Ӎ7�߸.�L=��Erڳw�u�n�O]m��˝?��]��#����߯o_ϝ>cN���=tp��/�.�c�����+W�g�X�ˊ���qXrq�.\�$odOC'yJ7�' R���p<���PM��3�ڀ6PIX\�Fqȉ���OT(��g3�4�,���쉓�6o�!�M�V�e���$2ae����jp�Ҋe�N�:�hɒt>W��M2ƅ�ق�����b�~�~����"���cc�"�������ɧ�@_w�6�'��>�pߏ��A�q"���'��A���$qeQx����E�#SGW����9+�^�fm����#�Z6d*��@B�pa�855�����d�A9ZR� J2L���2S7mdJ����[�d�C$�P,�0�U.<h�Nڦ,;48�P_�p�������Ql D���p[s[(������TUUzi����\zي��;/�	�^0aB�A�uf����/�w6��^���;���;o�!1/����՗h�Qg�)�4B�2��`9�@��s�d[E�A��PM���(����fp������� ��������ʊ���`8�嚫
��S�V�^?��I:;;�/���d�9���
�e�������/h��p�2�2����L�rY�@4Ú�ֆ`�[�[.�W,��q�����:w�#��]�fe8\=:<291�����ܺ�ώ��
�M�ԤL���]��뿹����ɿ��h���Mʠ��h:(r)[�9Fpƕ��m�79���Γ�K�$�"/I�AF�l� ��g��Ǻ���*����
�Tn��.DPcC���,�!��l��������Ň?q$	#C����S���Sk6�O �K&�,�Y�v�t4344�w�{ժ5����ީ�n�j�u{>�y�����7ã�Ɍ� 5^��8w>�/���S˱K��3���~�!�]"Oyy���| ��pN3��Y�)W#Z�,Jֱb,�Z}���7�p��Е�d��T'��l�gDr���%���O�fg�Gzfl¶��N��o�sp��>W��R� l>���V
����T"ɳ<�^\���WQQQYS������D��l �A��]�u�mnj���>uJ��%�g��l�r��{�� Ki�������m(O���;b�	���X��՜~��s/�M[dzA�I D��ǆ+"6�� �+V.��|ǹ\!E��4UQU�����R����2fa��s�$#{}7^1<8XUSU>���V��ɿ��#ps�5�	�b=��&U!_��j>�����H?����C�$�B��� ���)x3`��KdN�W�"+�?���O9�����	�3�<�`�`�4$�G 饱�9��8u2�M�>uD����c�[�\=;;Ӭ]����v���QB�/�L��`\�GF�<��.�����o��R|^ 	8��U��y$_eM���>���ˮ�ykQ�6�^����_f�EIwŊ���2�VU\��>���:::���V._���W^}���2�쏏=�]��kj�y���3��R>��2|m]}2�4I	��4���$��� %�� #B3��#H�X,�UMUmU�uDN����B>��yr ��0��d<>3��:���	���#�r�۲e����t]�t�����]�p���G�-Wm�b��ĸ�IʃVA5�mZ��;u�����O?�9�a�z�w��|A�����p��̰nR�H��y�]_<�ɑ�=�w�a*1�inh�䓽�7����dR������{I�yţ`�V���뚉�8+���n��5�VWEa^浵�fg�ĂŋJjqrl|�����޾K@(]Ӄ����I$�}��R AD�SН)���ra�B�����t2�phh$��2:>>RdX�rRgWW���8� @Π���-[p��%E2I�:� :N1����rق�j&����`Ų(��cGsK���N6uw����<����*�sZ���u$8��S�n�m����������oO>�@����؝wݹw�'��_5U#e\� I���\c����`I��8'eb�j�&٤E�ʖU��Q�H)��J�2�W*���34�/�O������C�3>��55��ޠ���F��ϟ[�|�@�pKK���(�&Ho8����ؿ͚���)��\���'&��*y��Oj�h�k�&�D�?��=�MU�m�>������9�١��˜d��W"�e�#>{衇�x�-�U�W_y���à��D!s��[���F+�@;\7~�J
�'�g��&,%��HD���@�?04�x������p8������ՖJE���㟘I�Ӳ��	J�!s<�AZN����N��)�@Y��SiN���[��Ύ��χ��������64֧R��g�www-_�n��~ �歛@W�"G��N�&�y�;w��<���@���/����M[.���~�٧���{o����h��wv���ƛ���E����#�k�7��Eΐx��^QՂW�&��e�\y`p��ڹ����~�Ǳ4F����Ll�XR�e����YM�&?�p%+��dlzjb�vmaz�SEF��ry��dˍ���Nqx���"O�  xx$~<�΀�7,_�~���uz�ίh_E�ERV.]625�"���tvt�!���Xk�U�~�[٫0�!e|t�ԑ�
r��x���^~�c��_{�H�����ɧw��$��TIɼ�m���WQ(T� ��-һ�i����m�$i��ǃ�A?���{���zN�/<�jK
拉�0A�w�'(r�6����45�P��A�%l�cGз*X�E��i#�s�4���w�J���z�[[[���:=5}�ò'�<�z�zZ����86>��)�T��"ҡ�$�w,��+6v^�04<̰��y�bZ��n���b}s����ǃ�=R�+���� 08��}�lwhx����!_L{/���HF-L�<�B���tfJ�����CΩT�*!%	W3KYrZ��y!�u�-�╪jz֩�P2=ɳ�V��R,gX�VHC�|D���c�l�W`>$��̻�������M�61>v�R��ظz�*���O?���.[Obow7K�����#�׮����ё�Nf&335l��Z�j��	[&-[�SW_'3���8C�l|I�ȗ+0���8�6�L� |M���|��y<iRR&>��'E������I\��Gz����QHC
�β!D&'gjk���d2)"���ғ��>����w�v(��h4�͖�%���ɉ12�J*��Q�l� �Q���I����p�ǎ��\}��OX��I'�n�����2LSC=�Gx^^�a��:ϷΙ��vI+�516<ف���ppzjֶI�	s㦍�^��5�޾�W^z	�$x<m�sY�Df���X4sɊ��.0J����"]d�>߆��O�:Q]U�`ޜ���٪�0v��~��[�}z*I��\��|�,7�������uu�+W�ܻ��h�"�j�`��2*�z�� �x�Bג%KQ �R� |�(`�r��-��9�A��++�o���Xʝ8uB��U���E��6����09=�L���H�'Μ�ʕB�0IT�e��O.������]<�T<��4��a��g�t���n���7�x��2���[k��W.Y
Y��C�Q�*QL-M-��ַ>����>[<v�8�1�L&���G?59u�8�8�dζ���;c�C���m���u]��i�����yttt�܅�,��� ^�j%�,�Į��W�Z]]S���*"��`��>Y2�D���0�r�$P�4�i�T'mb98#P��	�X%|������m^?/ȼkS5�����Tc34�b	����%63�ͤ����%}�E�ߴ�w�����!���}i��7P��y�B��{�QFN�f�n��;n�62��J_ �p\2��
���o@�޵s7���S�_}�e��^�|��MF���vc������"^�@f�)^*�C�%�E �����dhVV�trV/�I�cx�����{�
@`B���X�]�9��\2�MF���2�C�W*s���e��G�h�Z�2�f@�Z��O�nfڢ(k�`�77�������s����a����ڗ����+�2�r�|�u�\�y��hk��P��J�xE��J�����}����VUT4���w�#��O~�������z�����Cl9�����֪@�uMD�ɸ�K:9�m:�N��+{��b�X��"0N+�yQrtJϦ��B&M���r����J0�ñ�)Q���������&G2 �X��P�����
��P}>��H�.��k�j��Jg�ezHJ	�YK.�PŹF2�hiF*�'������p�_�8}�b�E�4�vF�HbSc��H�T�<�O�F�t����j�~��3�O�9�>�����ۻ��_�C���ҳ��/�R��h��v��m�،�kt�6-Z��/Q-,��M�D�<�� ��6B @�	˲�T��@��|y0#�-'�2�N�-�cb�/��f��p �K{|�b1��¾����͡\�)�� ���?RAzL%S/�{d܈�j;�<�2Q<r�$��������_֮mim�>;��;���M��\�҂m;���ڪV�<�$Ŧbo�x�&�jK�b�Axㅗ��$;?��0
�k�����YǼi�:����q�W�8����XSפ����PBNy��ܧ"��gxIr	7p��Iᇜ',+C�R�^$��|m˓��AFu���K���K�m�&/
�`M
�|3�����(��DBA*DI��$P"=4�����㏜�Ŋ�\�e]�mہßB`nڴ�wMOO?���LL�DB��=:1񵯴sH9���!�ՖQ�et%C*��%'��,C�w4������J�o�x٩3�S9W�
�u�� d��\�C�>\�EE6Q��ms,]%�>�pN��2�1W�7,0�#m��'�JM�=Q<�Y �d����'L��|۬e���Z��r4+aIK���Pn�P�m{���{�ts����~����L�ۃ�ώ����2��3�AE^ȥ��>�7\J�O8Bd,��!��3d�����M�%����T��6C��觀,��/ҳ3��&�'���Ϯ�|�HΊ��t�C�%r�H=��j���i��d̚L����Fq.$�K��	���<5eH�l�`*�q@�ʓ����>s���B�`+(S�"�,��6�Ӽ�KԘ[�"g��� v,X17ڲ`��2Ғe(A�~�gxt�"���$,!�o�e�$85�v�6��-m-�,Rb��X��cT]/���/](�5uHE�nK=M:�4;�^��_�Uj^���g�x�F�����OS�l0Mef��yUTdʱ|��Dp�fQ���&����R�e�ѶT~���r����2�;<hD�D�����֕��C�$�ƺ�m4K�A�
"B�i���@&��8�����9-��t߲%m#�B�f� �˔g�hvthttpXP8���4���<�"�S05�R���/�}W}}�����R��gG|��5Wo;r�pcc�ҥK_z�%Q �D����y)��F��F¡�'C�3�H��lE�����ў�.N���e��2��H1J�d(�=��ɬ���gӊ"M�� ��haX���i�B`l�%�N(�Wm�#��ؠ)�b�I��#<�B��e<Ju�K-�����n0���q��`׾���)2����W��җ���|���N�9�F�����K��TU^�p����Jq�&6lh_��8f���:x�X��9~���,ٴi#�8C#���VMu��u�1��m�8Z�����-��f��������H�D|&��`m�F3$2�����TZ7d^��uR��5US�lkm��'
y���g9�634�<%��:ыP߮%�T�D�K���~D$M�,�jN _��ꆗ��2xQTUݫ���d�T��P��&ff3�/�"���7l��2K�\��ĉ�heM�����i����	+���|�XYQ�y��o���e���>���gf��/O�1w~���]��J&[$�h��ӌa��.]+j���]Wm�P*&�G/������?�
!ˍ���AG��v�lJᅉ���׿��J���:��?�J��k}O���H��v���L�}����C�k5��Cӣ�Sw|��Ĉ�'��?���!1T�s����}������7��kǏv��/��$��k�^��K��A�y������Bv�E���^��+_~���rٱ��9���i@״�/38٣����;{.���=zPU��Hde��ώi�oں���}<���"�i�Y�����I�^w��H���-KAˇ�;gs�����|�k��EK�$�M͢o`�T!xc�c�?0�d*�[{c�cɀ/\=�֧3�d��S���.]0z�X]ۘw+�Wn��������D��[s��3^hk�˗���E\*9�{�6Z�{�-Z�d�U��-s��Q$ b�@&%A,U�ښj�ù�M2��*to����g��˗-�чgcSgΝKf7_�ES�B.6�'����]���嫮ܸ����'�Pd%�JE+*~���8�;��ϲl�پ�`{���+W@�ɖ�N����N�ڀ(Ȁ�X̾����nv�q&�.[}�,��x?�������Т������33_��F)P{��/<��օ��	�|��o�ÿ�;i��5��M��L�j��]���'���o~�����Զ�����K�wp����^�o�=p���7RӼhh�Ү��޾=�nN�B�_~y��`0��	b�;?��� ;�p��U�;~���Һ���.��Z�\_�̝ye�;+�\�Ѯa�����g;^x�L&'J��%��3�>�/��@��D�{?���ĴE�S���5����֎��S�����F����ohX�{�K�,ݻ�c�G�5��]�����/�c�׻x�
��_�`$N���W���X<�riE�h�tN�:�����|ޮ���7h���������853E�rۜ���ޮ�Q�f	��u�v~2��m9�������c����D��>�o�.XV^���N��W^|�U+�J���cP*�0Ϝ<�t���v>��?�ק�[��ʢ��eY�U@�,+�Q!AX�e�\�"_J������{﷑� ��gcj!�-�����(��P�iV3-�G?���#K���&2$�:����V����A�� d1���Ի���FF%�̇�4�̟�`ϧ�(r�)�.͙M$׭l�?!����2Z�qbuU-h��ډ1ȣ�:��3����Gr�TSK�`�����u�>�ܳ/��.�o��|>���82�,2���ݬ�Y�#B.��d��P���|�)���I+����|��|t�	���Wo޺�frxjxtx�҅�?���邨�ά�;}>ˊ�}�GS'ΜN�fu5oڑcG�v�'����v�F��� �z.v�?2��bO�M9�n_�jtx��o��sg��=�G-�9�q�.4m�|�E����S����f^��wu���"�#S�-� U���m���>ϸ�|A �������=c=ϐiq����A�9��llhL�AAZ�ʧ�9�=8d|�FB�W�>��p�b��K��UED�Jłj�6e����P��"� ���2�;�?��8`�bhIP~��_��=�}�ȁ����y�X����GeYJ��^���%��(O�;^�����f���@������(H�t:Xy���w��æXQ&�q|�A2e�pH����w@�e�$�~"~�L�Q���Ϧ�0q"/�U(_�gK}a�TCf]�LsXN��x�`����IӸTҮ����8����K/B$�������v��v��� e?���P�#C�bV _R�#r�}��W�y��;���u��qv�� �'r��(���������ևgv�v�f˒�,��n�ml���Cυ4��?ܐH$Ԅ�L�1�w�Y�$�ȶz��>;�S�s�1���Kliw�}OyN{�����"[��)^OBǎH��(�^ ����؞��0�1�[��$�Kt� �-�b�B��q���tL�cϘ.HR,8�ҥ��~�d$8�"p����|#=�g�u}��9s�϶�ƨ����23u��o�%3�s�䱝��j���̚5g��U�pB�����cr����"7e�䂂������ԝ;w���z�����|X�3x�@ (�]�a0�O Q��#����$]�rc�����9�^Ul
k��FBK��,M�il����c�#j$������0}�H� ��iҫĂ�`�;k;�BÅsj,hï��v0X�&�|��&�͝�`�4OR��+{~�9&wl��N5,�3��!V d����t����hF}���h ���7��^������6�I�������h,��?�t8웿ڼg�O8Zc�d��xH�vd�����C���9Pd&�� ��uL�`)L��ck�����/c&��f��	�$D���Wy�L�P��
��~`"���">|��5�b��S��H�7v��m�y�O&�PYQ�	%��������L�:+�(�F9�Yŕ�p��7��={�f�&_�a}WGW$�D{rjj��\iل;o����;C��A�q%+3��7
��Ǝɶ:|1�`C&j<��|.1�� 8�ag�Hr��*�S��:#��	���D�(�$D*���#Ϻf��8sG))R�'3�5� r6B�m?b�fcCa9?�(�9q4����'	�d_Q{�����Ӓ%��/��>�7�Js�7͛�]�;c��יӧ�RRW�Z9k��p(����3deʔi�,]Vs��p�x�b��z,������)+qB��ho��;!�qQt =7)���}�&\�:)<��xdd�A�0�sG@���ԃ"��I�a-��Ǧ����ې����whR�׮:uBs`���X��O3c�&wl��F�_h4�P
���p,�S�؆�Eo�t�ʵKϝ:3i��vlHJ��������𸦲p�˕>t��������B��3�/����x���Cn�%�Ր���?���7��D5���q5Fmvw:zl�#v
M�WR�1���|�8Bg��,*o�bȔ&�y�! ���H��s���_�aK6E`E��}'�	�Ȕ�6rL�e
���e%�ڱ����W�Q��!Y�d�9	�V�;wo;Z���b����w��PoWg�����ӻ���x��n�����N�&784����q�5���a�G��[y��۳H�v�=(r$?\47�K�?W��3�q���`ӲU6�Va��a�V��&�xV6PFR�'U��'gNS�/�Љ���;�$6A��'��h#ND�b� ����p?s朙3���B�&��w;�M�ʫ�$�������Z�x	�E�GF�l���x�FJLg��|�1~��|���(R"&,!<1���A������s�PZBS�` �72�u%W�}��W`Ll���l�IFzɕ[�xl�6	U>�YA��ђ)]@J?�p%$���H����xt�i���q�<+�<5���.�0[�'����&>�?���r<.��r�x����p��
HO	��ˊ�a�\<K��S�%h��Q@K���L�3�< |�I��9Nd9>�DAL�8C��&q<�s����d�g�R�MM�Ig�ӱ}ݒ-�q��n�Z�wa�E���=)
O�F¦X��*\W����@�݉�,g#�la0'Gb����U��s$�^��Y���V4mp��
ރ�8�z d!ё|����A�߷���Mpp�S'�X� Tg[Ǿ}{�9������<^Y��ƛ���?Մ1����C�v���###cƎ�%&��.������t��urV9��4C�uA��b1���e1��I3Ξ����y���U�y��v��k`-,Я�
�JʬKBQ 3
"��ձ}�֡����ًW��6�lBW�d2@����A���@�&M(�v�������UU'��ǀ�%R2�W]���1J$�b����yo��O�����/\�dio�u_p�����G��2FF���`���$�=���������|�4�ı\�T�!�Ҵ��|�S�z8�����i�W1aaA��U���1lL�i��H�A"T��@���(h6b_HK���؁��w��V3���YM��X)�)֠͌��@0�������K7^�8v̺W����=������H�������\�����y��]��Www��۾e��MII��^򺝱h(��:��=�++��1��z`,;e���D�--CZ,JĂ���q�2�O��3�� �	��U�e(r$u����HEh2���~�g��C�!��c��p�u͗/�'p�I�i��u5�{��p4�X��66^:��g�;}����~�(����L
�.Yr��p��}N�7�!@�����vV���^c%G7/Y2.ol��1 U��z��r�Ȉo��2���#������WRX����`ɓ�������D2�C�W�	e�SpP����HZGآt�m��E�Ȉ���F��-�p4�t:U�-xq��X���[C T@3�Q�"q3'{\NJ�M<���9�����,���ח_~�w�Ϟ�u�E��_F��.��r�i.�.+
R���e��-.-*N�x~��ӊ��#���i)��^vv6u!OK���^n���H,������y���瘫����i�mpc����UKL�̫�B�Rt��ìI�g ��Y��j��B|������8V�1��b������(���Ϻ���xfd���q�^r�n��8`N��mk�p�1����=�d�JOjRanf���ٗ{8z�	�۸۷���def^������r{�.��w�JKOj�肘�>&J��?�(	|��Fe�KN �@�r��L	��$�k@Ǒ2�]E�@�g�F̙Ih�����ȅ ���(�i�I���2~�td��ppZ����ޠ����@��f"��z<�p�G��x�D�?�rJq9&��d��AÍ�odh����!6)��?�[o��������u맲�=`�Ξ?K7H�S� 
Ý���f����Uehx��E#d���2`J*>.���*�m�e���lH@��:���bG2Y�*�	<F>���K�r"E�6�ou�G�id.>Y���Ѳ��8��HTtH,�EBa�_t"�"����E��2�N�'b�=����p]�}���Â*S J9P$;Б�ٓ�Ȱ��c�L*A���4�����ǎ�>!�$M�1��6�y��
F�p� A,���4�b��nAj�b��b+�bM���2?r\B��	��ߐy Y�L��ĳ3,aC��p���]�#�	.	0��pM�W}5��;A6��mf8OK�H�.:=5PK����[�7�H�Y�(�V�8�L�]U$�~���2�i��.j���9&�"'V�)K�.��%Ό��=ݟ��1�Pdӭ��M�(�`�l���nٲh�������~�i����=���v�ei8�"�O�����7�L���.���9�������?јL� $U���� �'"
Be�BDk�Ȧd�hӲ����SzLP��7�M�y�H~G8d�k���u�M�,c�#�raQ�}�ݛ��R^yl��ݠ�rL�7���ZpҒh���x�\?^.�������{�B!7���e+�;�j�������.E��ŉF�%�gg����"���"$��G4kni�	��0��6� ��%aB��Hr{y��=����)i��}��A;����:(�N��Vz�ęVo��ě8bI��h�����/��x�<�����x^��Ukָ]܉���_|�Fb�̜���Z(������S�z�ч~xђŇ���ƛ~��_���ر�xOU��3��>s��;n�G"�EE��s����Ϟ;3m�Զ��6n '����>��'�Z�]N�s�>�q{{uc��䔖֖���J""�Ƒ>�Faz�U�D
̸���ٰG�%��,6�:��`����F)xV� ���oCr,�X9$�e5E]�lEII�@��;��ڼ�)+֬r'{͘�i�ʗ_�k$�gA��&������y=����r�M�~����:���s��l�~+C�L `9���@U�-�ӓ�$� q������ʹ�7�_���<k�LM�D#����vI���7|T(�GR�S����6�c�����*a1�qE�.�QP��6�ue9N��c�=F���v8%���\p4#���1��/�9��	���Š	����˼�ʫ�)ޢ����k���ם=�d�������ρ/�[�2�[.G�ص+V��'zq�ԙs*+�V�ZfZ.
!#	��h���0�P��>��Fa$�K�����'d�����@���#yy+E�0��0�yR;b���T���&�KLO��������DS{�G Cw���� �c2�����m�����O�4���H(H������Ug��k6��_]S2
�x��߃@tuw���P V3Fpo JIIJNr T%���~Ҕ�p�������_�#TS�N�eӭg/^�}�d��P��z���ٽ%�'�%�����<}dd����)��x,d�0S��Ȳ��sg@�/\:�=~\AWw/ ����SY&�DQ�8E�A̧�W���#G��J�R�"��k�֪��ۙ:eҤ��6+���ڵg�k��hb&q*Y�����nݔ�0��w��p�!�E5yÍ�oܰ~x`��M��_=u��bꌩ���G1�d�PY�d�A$�ꋯV�Zy�����~���2��o�ۚ�����/��@ �)�jG"b��"�u�^�s�$Ό���4����Zm/�p'�6k���^V��@���۷}���� �c��C �˨��6�3�4�\4�2y�]w�E��~�񸖖��*��Ə?�fּ醑 ��T( �]�=��5��y�����������&O��"++��dpn�ݮ4_��������g�����xn��%�iۿ�򛭇W�]�9?@e r[��b@���8�3A�E��7����!�����p:��l�M��\�6����lL�$9@��3Q�39������8	�r��_>�8�_��-q��G�!.�2���)�`)´e1��IPy}����}x�19Y����R��Y��p�f��p�T��NIP�8�ڴ��S�4s������i��V@@HSy���p>FŚ�jI��s:����y^���%��i:]�pƖ�5���$l�`24B���</ja^2��H�.+'��G+�gډ��X;�Ñ��J]��	���C�������d�rgN�!w�"��!��!a�����[9
L��Cxb�j뱙��5k&����hX�U��u�E	 d3��&��#֍��I_��?Uj��Y����fPK$b�a53GX��= �8�$����kv��.a�*n�aF>{*.� � �"}��5&��m�P���1���@�0I��˱����gO�
BE��+���:�S�jgG�����H4�]nIC*.����3.���rDg(2�)(̜#S���U2<"�j6k�U��xʸ�D�$  %'�J�Tx�X\�x�����H��;z�`wG��˗���V�Z7vl:@�ܱ�|����cJ���3�Ы�-�H2,�<%�6A��6�UNO��x��.�����x�X��@)"��(I��U��&��Hy�޾�n@�*AQA�`���%�Mq9�OE�m���w�}�7)%��	�}#/����?�ݞp�@�R+?���U��E1��ޜ"�����ra#��9�EP���'���(}��G�=I)���c�����?����4)6|@8�d��)}ݝ����/M�8iLNƥC>�38��q�_��<e�*�7���{o���-��Y��w����X0AGG�{��;�}�j�� p���'��M��4�4���8p��h(\^q$
~�E[vf���e�G���v������ޜG�4!����";\Q���9>���5)q0P�->+2�YQ���20\�ю���1�3q� �:9$���[�ch�ᄐ%���b�xhh85�g�/�v�ƍ�`x��呀�/���pL�9+{����>���|�7�cC��¹�y��8B�Q���ܵk���8���������$IɄ0H�K #o�!w�8�R�RO�:}�ẍ́�IǪ*7^����D��pTWW�,�i�X�/�����Yw��2�Y�'��1c=n��D�F�pe�ך$7�kl��O�x=(q`�(�J�`g1�q%��"�61Ws�?�u�H/iQ��p6�!��`o8�n+������7����v�������������H˺���+��q-�~�ңA ����4Z�3�;o��h��-�~7<��p9��Z�"�����Y��ڣG�X�!N�=��gd�N�/�\�7�������c�qLo���p((�cH�(�:����$��EeD �,_x�F�#�J��%c1�iA�L��=�&��r5����8[0S��H�gX �`�a��Kf�%�fpw���SO=�� �K (�C��yY�cM���Lal],x�sg�/\���=�lJFF��E�pL��j�ڍ7���?�����`86��������h��)8�n�g��Ξ��/��+� ����z�o�i.��ps���I-W��pMm-�̬�̃{�Ƀ#����p���@vR*1�aJ�6 ܋�lb0}�1L��(�������2Z���۴p8���4q�ԧ�|��O?���u�w���w�l^4{����o߹m��s'O�H�_��V�X�j�@`dLN�3�������q�w;\u������Z�E�����_�|�K�핿�ٵ9���I�'�_��x�V�n9 q�4�3&;%%�W�p<�bЂP�vq���kV2�^�-,(��k��ÏhME���7�de�\l����!��r,�󤽊l�68�M�Q�]�UO%�l����ix(%$���p���឴����	�&��>u��O>����͛;�����$CA6+��P��ΎÇZ�x	�(����ٹv�Y���������%+�eq�K�_����_��#7+	�#� ����Ap��Q���=�F�� ����;��N#�;���Yz���qMknm��{#8�$�&�F���޾��'�~I��Ѵ Yp��������pJ��&�)"�*��l�2�: �n��$�&��4��04�!����))-�H�X�h1�r~~(Dv��ɞ�����W�D�q�����V��?}�·���/������[���k��/�SXU��v'n���_Y3g���� OH(9S;�F]t8@#��gge�t��������{�h]�m����$�����d2:/`B �Gҡ��&q�mVy$7'�CS�XS 0��W��W��f7�8i �5צi�����>��ȑ#�gͪ���<~RÒZD�j�x����h	�J��������A��Vq��@�H��� � S5�U�Yy�9�R�q��Eʙ$eG��Pm���^tHԳ��cZJ��x�÷>@"H]��8�?���WB�ᓝ.WYY�}w?`�ӌ��QUQ��ޑ��~p��|h��L� ���yֱV�q����~yt��ekW�v8��$O4�p�2��I"/��piY٧�}�rzFA�w<��>��3�����=e�L�!$���f�H��fuN��u�]8�L�<D����,.RSNd�͛㰋/\�k����-�t�b�\r�1�l�%krl��v���.��^o8ݽcgy�����yZA ��鴧��.8��ޮ���^�����3&G-^t�¹��>�œ�(��u3��M�@1W� §�Ϝ:c��p�
�p$3+�`{G�,+����%/6�_�va���D"a���t���xiٔ���&�PZ-X��%�H����2��nv��3����V��3O?=� <�a�?��s��������bٔ���|���N����9$\�?��cx>� %Ɩ-���kVH.��8+ٓ\^o����G�������ʬY�ep��'#-�u�~�ek �+�K��C"1��PlH%�+� ����'�<~�%���t���p���`�*{:Mwv������ƭ�2&y��*qٔ�8NE3T�ǣ#5	fSոJzu��������.X��h|v"���o�؀�-Y�4{LN[k+��N���C?[YYy��vǞ]~���t�%�IC�^8b@᫖-���U�OGm�����x	�r6 Y���pL�8F�=�����A2Z�{Ig���lϷ�)�ɠ$�` �����]C�f�T)е_w����6�B���Ʀ��q�����ת�"o,{�$���DC��,�̍�$NVyZ���*`���+).��I�;v�3cfBQ�o��?�7U�dIk4�����)�dP�ۍ�VM�ď����L()Y#Y]�j�����6uRIQ�Ž�BƘy�<|xמc5���z�闚�bJ"+-���s┉�i�8|ENN�����pHQ�bԾ{�O#�>�k���!�����
)���AQ��;;�����'��6����j"op��k�G��h�,�m��V�&�]7I!!=�	^t]�}���ֶ@x�n���Ã�v>i��Y���w���
[��g�9z�ln�[6m:v� Vzmܴi�J
�O�k��˯�����$�G*+��_|A+a��ԵF|i��9�I�$��"����@0 �q�W(���K4����3N��;:�~����x0
���R��{��0ecb�EG����J4,�Yt�8*�2�hmu��ύWۀQ��fP�Hj�6H�����dy�� ������~�ػ ܕ+Mc�x�ۇv�ڽi�����l����Ѯ�vMvF6��o��&x|��������M�ߺy�fxĄ�g��%_hl����v	�I
�Un���$�чpg�w�q��Y�|��{�Y�~4�����i�-ޠ@���T)-�D��8�\�a u[4�X�� �`_���H2��=I�]4��A�
)u��:��|I�)��2�8�"	B�4�Є���
v��7^:����,��ǫ�o�mݣ�?<gƔ�κO>�\:i)�u����ʓU���Ƣ*A��8������b��L�� Dn|��.����#4
���󍆂�-�/(�� ������.%��ǎ���1�� L`iF�:v�s����zA�!`���x�P�UkD�`.\N��C�C�!��!(ƀ�q�C��UM��	ʰ����b�j"�]8bl�čz�i\=*8)�G��y�p=�H���g���+��vGGw8���,�"�����x\���$eNPD&���.��ƥ����@�c@s�j����5�.ڥ����ӧM,)�[��?c�b�FW#��7_�)D��stk�!���MJR�q]U|h�	P�(����	"�K8����$����i�x)%�#'��.IP�jFv�[�C�#�j$"�ޠ8��s�xs�Q���6��I��k��ٳ�����Dў0cH�CV0�'�d9Fì1���n�cxp�ȑà�:ik�-�&֖@���IL�aI��NOO_�j��m[����;��L���n���o��,	v8�;�)�ѩ�))�IC�.Q�R�5�Մ*" ���쾁~������ ��{�L���}ý=��l߹��x´Ie��5/NA�-���p�$o�&���͐������d58[�;<ĹX�5@m��o$*��H�
Y6���n��x���1�G~���mʴi�(lݲU@�,�h��p7y��.�i1��S�?Y{��9I��9:����b�G��E��{���{��}׮XƐ������=� �PT��A�\޴���L�z���E���TO�>��ܜ���cǏ��uwє��#�-^�j��m�O�X��C��ò�i����ҷ �RpS�f����p�c�ġ��=`���$�����uh��=��*	��r>���e�e�����! Џ>��[MKM���Oo�n�I��`����>`Mo�tkwwgוv��I$���ݺiS]]-gL2:�c�H�@=Q9`�b$0)�d�Ý����w[D��������Y��v���|�FqlsG�ȹ��E�����6IA(>��˟�큘���C�'�{���L�C
�}C!o��nX<�C���yXX�:f
���0py$`�;����Kv9�^x�/��l\�̙��������V�\��cUT�|��w` //�λ�;y��YF /
Ԍy���3g�f�C����b���L�:p`G�EgʶCup��#�4����'	t��i�S�S��ɀ��t5��d���q�9���Ԝ��� n�lik�rINJNj��Rx(�������N�+��w&���"�㨟HS���ܳ��ǽw���ί_�6=9����歹��]��m!�Q�  Z�;g���������B8���¢P�#����� �m�w��"�Tw�~��΃ TW� �%���� �7\}iQA��&瘽`im��3�ڣ���6�$�UU�:��':Sy��.��hk��DZg��Bw�`�n7�c�R���w�QVX���s�E�W.y�����a�k���2�5\�Bf�h��K0��Wڼڭ��֯[7o�<����?��E��m�mz<1q�T^�̜9�ʕc,���$�7�[^^>nL��S@���}�ɋ�,���;y���s ����}��922q��S�=�����ȉ�g̒�`ZJJ^��`���=��& 8F�#TV ���`�?z`���)֢tL�P���.���(YG�O6������9S���_��w��yN��SPX ���������_��SJ�N	�	�ʎ�q0��M�Bp�����z���Y�gϜ9c��@m�WT��N ��.�g�������u��.)++���������'j�XV9}�������8w�[�M�p,MMM��`�YjVs{_AaQ\I���5n��w>ٹ���͈��8�*�Y%�b��y��a����5�%-����m��Ge�@�\t2��Si�0LwW�'�~Q1��JJ����˕��}���+���C�N����������L\������s��ʚ��c������?�:�ǆ�s���(��}}`"���]���5�0?����mcs���I������5�,�t���C���k0�J^��㋋
0ݦip�&.``x�����<i
tWW{j�X�h��w�#9�:f8߈��88h_0h����T<
5A�Sٙ��͋C�X�QH����.�^�����l��::z����frrƴ�E'��{{c��z�Z�dw4��%;3�RsKvV�o�y͒%pu'O?s�'`W�2kV�IOK+?z������?�t8��Ql���h,�$�R3�i������oN�:)/;���+�.w��ƭ. DA���ٳ��Cu91�O�UU�/���r<����GZn�I�:]��'OIa~���HԎ<\�g�Z��ҋIn���HL����;��g_���F��KD�T��d9	 �]p�\N�/�Yl�)���dd�������C����Ǖ����׿Ece��C�k2�h���^ 7x����q9�/a�9���=�Xnv�؞��EK�=z��bX�ưt�.9b�0Ȼ�d�e��JS���pi&i\R4�!�	׾��P�/�����;|8��q���q ,
c*�]w�������a���.��o����'��v� c���IKrA��v��u�T�{h#%A#ɓ$�\����i��Hh\o$�!��1,���P6�P)���-fge	� Q�!:~$ڲY�R.	�#O�����o����5m��5��z����o����=67w�ٓ'M����%;�!���H$���d�글Q'�XcI�������!��%9�=Ս&n��RV[lQ���	MO(.9U_��>#�h�,\P]U�eIKK{���"�t������5o�r�,�����Iz�H�"e,3�]d�=	d�\���vFb*��C;L:���ⲵu�� ā	�%I+Z<
 R��9���18S�),.�O�ajG���'O�o�b��#�xA���l@bbq��k$��d�����΂��2����{o��e�Sg�z�߲K��v��u�5��8iok%['P����f�HB&�w���n�+HaBvj`@�Ư�v}��q��1�����X��mP˿����J����̜�@�	ql���Z3� r�R4?4샛��
�B.^�0�p�?W�5pdq5�,.��^�p�'��ţ���F�U�{euE��: !)i#C��HX��)�IPF+8C��4���U���O?^]��?����̝{�M7��C��f�j�����+q9��<1sZ٤��O45]Y��	� �`]"��O�'�S�r8 �p��q}������X�����k���������sQ���s�rD�>TC E�81�ێ%!�E�
�����"�r��.[z��
�p�L����+�&IM�d ���ͻp�Q�D�X�?ġ@5ΐ�v`d��Iz�OL�,q��Y�f%��1c�=v��u7d�$�ٻw��w�yG,����"eqQ���KJ��d�ɱج93���`Hٽkߙ3'��t�?2�5�<N|b&���Ï?F��qw'�����dtW����v���;�n'��od䮻�
F32�c�� �(=Z�p�6Z��ݠ�Z�0� K
�PN��$o��� i	���xL޹k����8�C�>���.�Qd]0���d�X�ˮ�ĵ	K���q�#kXSb	͘;on8ܴiSff��#�fϜ_Us�n��1e�ⅽ}�&FC�H���tϞ9���w`��t��c�@ Na���u'�D�ӡ X�Ħ���rs�ܵ]��NQ\�t݁�GX^�q񘑜�r��
����>8���sr�xB��G��t�"����j#���!���m���@����p͋N�0�J${Rf̘p�����L�H\ڊ݈ۢ�T�MJvˑE��qZM�"gH1��]��d%�Ȱ1�Ht���W�'���o��5��2�����Ӟ����R]q������ 4������,��Θ�`ќ��T lՕ�XC4t�[ɠ��nI�׮\��+��7��a�X�b�_��ē�36+㭷ޱ������jkN�_��@��"�;ְ!�5FY	?�=�@����3���|��+��<�g��UWOg4+_08489;�$��������X<~�Թ[n���;�̟��r��g���f!A����=d�7�m�6��������􉅓\�o7;Y,v�+�G}<{��3BÙ��@��I��R^Y����ookK{� �dX�����a��q� �����'����}���5#�Y�P ���I�>��D�R�-_��:U�x2^q�=YGq�)�):k�*�y\w���2}J�ً����Z�.^c��L�1S�m'k����)ӧ��q���$88?/ؗ-_�r�{w�ɓְ_zi�ԉȶ���p��D08f�P�����U�|��5�Ϝ]��B�
 E3�����j],U�����S�����p���c��?���Xm��}�m8�Ec�u���hX����n�-�o�����O(������t0���o�IMF�?�+I�I@�6ԉdQ�a
�H�F����v��IR���h��E���9z���l��k{�1Bjii��i\w7y��1cs"��쮭��ɒBp53'O�fmW;%�\�J�[Z�:�>�t��I`Бגt�M�h�Ý�H)��l(��f%	N3A�5�m��a�=������)â	�o�!ċi����ёy��h82&W��0�)Oʊ���ݵ�C�"ü�2J*�d��HvO��H؀[����qE�����_����uUG�1��kb#q,x���"7��f22ό��u��#�8|,�W�'��L´�<�8˘6>���<��e\�,򦦁^�XS�TY�1�!]�H|L��+�>�1g������+��b1�W:CXS�]��������; �'��e��g/���P�b�\�dVl{�$IPT;�Y�W bƵ:�]�!Z���JRO����)	B4;���k�'kL=���~�2)5}ujv"fD��"'�"����Gx �o4�����d�Ez4F�2�jY�tX��{!M;6�)�J. Fb��s\�aCzJ�Ç~����`���暴�T���u�-�d���)�!�X�ܱswgWϴ��X�x� �z=�@0x��$�I��Z{�S�A�����<�h`媕ƃ@����\:���|�5����o���`��3��**��^��aw��A��>��n�ycF�������؃w<R�b��c�=�,��U`I���!���`�ˆ��6�t���Db�G~���|eM5��u�����_�ӡ�w|��!��K������+M9YY���f8j��]NG2 �>����`�ҥ�>�"	"���B�W�)���kkk�z�fϚ�pѼ�G�S��"��'�<?5q��`p4K̛7I�~f�q���	H�=^8�fձj0�N�,{��y��i��H����UY�o�~�Ӧ������]�nݶ�;F�?�E�KÐ���\7c�@\A�q9��P5�$k֮��ˇ�\�l��33f̸�����
�M���L����hlƬ�O�PBڰ�o�}Ǯ=pɗ/]���{����'��̼�> o?���RS����-�B�iJ�FC(����V.[��ނ�T¡�$���={�[o�)H�HP-�a,�iȀ�N;�:1L4��<I�Z�@�I$�~+#33��tG#
����~���.�8����l}m8��L�'�����%p�r̴x����u|0;8fA:��/_i*(n'%)trŪgඦL����o����ɀ�1c44J�r)Y!S� ��h���?�DI����?Nd�c�g�yΓ����׷ݺ�O?+-�*+
��z�DBy��W�?�<0��ҪF�6 &�F|��M38BFb#!f̞)
B���f+��t�J@�ǫj �T�x^޸윬�� k�7JǕ�`������Te�����A��`�"�p0����wϟ7��h�7����H���5-=5yph��d��7����ߓ�(�ؓ+W���}Q(--�x�bB��~ ���#)I�w� {��c��G�Q{��j�?���Qz���cr�tuv��_��#�i2��?����a��?Z:qD3 �Y����P���༫��;����x��J>���v;��_����l�;N7����wy�1�e�^d&)%M�5�A����'M�|��(�*�8<�;�p��?^�%+�y�Q��An�;ڝ.��s�2�<yʔ����E�{z::�/�7<����f��ğ`8l��u6n��BCäɓ�l۶u�����7�.���qP�v�ex7��@O�[�-[�ldp��_|t����҈m��?���._~͎;x�v�J�`펰[�]����g����aN��|0��d���8�p$I�;Y���a1adX`]�EV���O	��	G�7_�|��e����E����rssrJ�oy�A��C���2��\` ~�X\���l��9E�!Dq�^����~����+���w��C;~ܹ`ޜ�{�HX �d;s�4׹s�,�ް��}۶6�_	��?�gϑ%�7�Ձ
���~��g D6tg�+���ԟ�x��H�0��CZ�J��C������9QU^6�L �����~l�Xհ���Ĳ�k�#����}�p:�b�v&a�@2 �E�%gN�saʴ��NTT��o��s�g�~�c(�Vn���T""��a1\щ>OIh~����`�޽�!�������G~��_�<yrxx0��{��_o���V���~ߓ�m8�.�n�]����I�j����L |��+OyLb1�$�9��IR��U�2����{(���:�^5Q[{��Ԋ�cֵ�'��+Z�ryWo��'�X��t��u�0��ό��(�
�,�\��а�Fw���&n�����T���e�``}��+�h�A=�^���󏂿��/���%�8��G�$���՞�C�$y�}�Y����"��pQ��ݒDe=&��\�!?��q`e�+	͉	V>�|4a)�y=��E0�'8uʔp(��m^8銊
,GJ'��3y�d��.I��.\8����E�u��q\�M>��,����64p��!$��WW����á(���.�֝L$@��A.��[<h�_�>mּy�|#�v������wߵ��;��9���55.%"�ఎ9" �L8�H��0�K��.NP��ql���1%�׉- Z\���f���ʊ�֎V����iS����@s�����vs&8��f͙��?���e�Ν�x�q [����	Ÿ.��Jc,�G��~��ჇUM!13m��	A?	 � =47����r<;+;����8	�mhg$�D��vG��'�	Lp�2"�t`oqa~sS#/:gL��p�� �q%>y���?�l$4������5�h�)���Dㄏ
��$�c\n.��eK?����9s�\�~��g ��������~�e�H8E�/~���{�����č7ݸ�������%W���$K�e����}IN;����% ^�P3ajE�	@�tB�����?�#��Dc�����D��m��p��
�}. %�q�p��+��T��Ǖt� �~���Up�W�G����������?��Ŕ̬����-_�t�T�M�Ai@�̰�@��M��5i�$'�s�C1�-ľE�n� ���5�ӦL�XML�6����t=��p��5/��wX:��|�J0胃��>���>^��ǁ�_x��O�l$��B9����^gFZ�1�=ظ�B^֐�p:�1�2��V8.������"��v;�QN� �p6��J
�;�ZEkp�E�/ɲ'm��y��Ԝѫ`�DWW���6��9y�
0h�$���h�
��/�xs	8M#��a������Db>�0�FB����v45����9���ڴ��*�pKτ�R�2�G��rζs��̴��3g{�bc�o�e������/��7�1;Bg��a��x��%T-j�lO{�>��q�ڵ�=p���ڸa���~Mt�����#���`y!
%'%G�QL���k��G�am��S�,F#�������V�u��8����qڀ���<n4��p9��G�����~�b�� c*Ѩ
�kC>Y�	+rb|��e˖F�x��^�;H%Xl����k��>%��+�BՉ��5�=��\ʢ`1/��,Y����97w��>��3�B�<efLƋ
|��=���q����6�-]�"}��kxNH�&���Ia�Ý�l��R^z�O��]�fqA�ÿ��/{�M\�3g�����ּ�#}}pr��M=u�vɒ5W�4M�X�2zo_{Gx-��+�.����[Z�+qu���J8���o��PR����:��ܕ�D��x��W�mnm�=��3D��Ȇ#�+VO()ݻgGk����gtww��5�{�} ���'�����)󜨮ƍAz��|���n�!ɕ��G<z�.J��a%[�|i8ܽc'�s���3�J�JK�����?� G������{�s�:�SS���?���\w�R�������Ј"{�B=�y45^\T�~����ݽ�~�=�����G{�֛o��>u��3�������ҋ/=��/o��d�TUY�������N��.5�KO˔�|^n��)��"[���c�OO$���lБ5��������SS�a4q`���'�{��̞�%���7����|Ѣ���n��;ޤNVTd$��u�$R[�����=�ȂIv��U�����K�8V�6o�
w��,����3lŉ
���i�7�(���z�'U���ѡ��6OR��D������J'&�|J"���dp�I^g��9+V���ۯ����?������0�pg��بZ_{��R�/���/6,Y8k��ǚ��D^��jvF��?���&+2�(��z��R��s��4��DeUENV:��KG��J�"I^o`�wpp��`�#"�5��z�ʥ��0 �v�ڞ]��?X'.k��R�8Y���v���h��@�B����bB0���,`�����$��p 'mp	2���hB�S�m,x}9�����߿񦍡�Cs�o������Ec�͐�u����H��q��-`$������¤xE��<%�J���7l�`O��B8e&ԁ��d{F"�����3v�7��Z�jyY���{�kjj�Θ�����������i �����j�!$t���E֊} ��������fyr
:� �PB�
��jjiI�Y3.�\�,�E	��XsἹSJ��P8g��NB�db�IeӪ��A�9���O�D�Fq�h�����/(,���6��QÀ:eY��Er�����0�����6�G6�	S__���~ ���C�$L�������w�o5l���� bG:�[��@���sJ�H?��.!�Y�	D �����v�
L�T � cۚ]�[\� ��2@uPG���8�Na�[�<ix�σdR4���v�w|�u��ukTVVR�-8N�KR2ec�/_i�m��P\���,GA·�qߞ�t<8�,�c��nPo��-@��e��B�`Ч36wr�]J�a���n��p�0��a�h�)�0>�����zd8)%Y�i��F�pf�$�i珻}��;UD�hǱ&�(���8u��2hޠ���Á +1ӧLf�Ho�@<��q䈽võ"��e�#Q0yY9Y׮]c�͖�˽���#Q��'���0=�a�3�<�D�N@����rvfm�N6l���hwn�q���]^�͍Wz#!�k�<N��}�` ��!t�c$�7<�6I��*��7WCG�+'�߫o��ϛ�w�޸��N̫=w��[ow{$orJ�@�̹���Z38*co��BdK1�I3	5NZ���c<��"���)��:ޑbs%A��p���8"*HM�V�ɧ~�j�ʦ��3f�x饗S�����C�TT\���>��0��e˗�����.�/.��������!�'=�W_�3n�g��E��8�N��y��Q�M� NsK����B�D�F5�|��*,��*1�c���Ĕ�%�0�����*)(P�A�S��<*qt[c��pB0�ȑ��|�B80:q�1�i��N�3S3�h�!8��:��@A(��t�����,�qrX�5� �Ǳ�?��g��i���o��`���{B٤������'�|=uέZZ2{��ݳ��q$�x= �V�Z����I�^�iȲ��g_���2����6��F������MJ�(�ڀ@&TȜU$!�a����c�`R���LJN��m����ZU��]�F��j44�.-�ť� } )n��!E�����q��C�͠:�[��f���K�H�qF��� �=ۮ�TR�DI���w�đt,a����?Λ?@����qx�:��,O�9�aO�$۵8���M�MKW,����:�/���������� 	�������5�o0)�3��g��������%A������7;M��Yi!J��,��x��<�ӡ`�dJY�9	�RSSC�H<�(�8�P���X4u$�\n�,Ác�d�5��
aE'Ɏ���+�������=��$d7	&$A B$ �W����:
^����vtj��bA:�juF���#Q��" d �#��;�c��}����Lfgw����������>R�D�ɉ�&r����7N����Ƞ� ��pW!B�L3M��G�ٿw�����k�X��+Ǐ�0�-A?7�;�!^n?��62��nn.����+��=rd߾/XQ/{K]�To�/w'��uM�mf��k_ў�"�'�^eyil�p�I!c0�I�3ҰE(�9/}>H�M�����Na~(�L�� 
�Ek�Y��Q�cb:��X���x�y��Qx��� ��_`�6�G�u��4Mʴ�f��� @Y�E���&����A�up��i��T���H��G����EYT<q|��ﮟw&
d��}�|�?��2�'�u<ɴ�u^y�ϯ>�����ä�O�x�sH�F��j�x�uy�����TU9�FwMdlr\ҤB�����T�Ʌ�������20��"���X*A��iJ���'�
C����t�>�kh���&�~F���q0�"R9�JѺnV�<���+��)"����h�~v�7GOv�����fΨu�T
�x����=�i��H8Da����?N����'����`����	b ��a�o�Y�;_6UA__o��7�������G��B� Ȓ���K�x�B�;F5��h��|�$ˤ��;H��9c|��]w��u�񱣣c�(���j"�B�d@<GNb ��cJ��uo��� �c�����x�P��5YZ�9>���ζ��Y�Ș)=�ϭ�^[UN0OZ6�/c�VP��"����s��R��i�ͺt�(��3Avu}���E�4p.�홐9����Ւ�P���t�ҏ��r�����H
4g�AK�6�����W�6!����	�$oX�Zi4�g�><J�J&Ƒ���$^�B!$��Ei�~#ܼ �R(ΪC��}��˰�l���-�'�Ve=��,<m[X	B$�,s�a|y�����P��4��h;��"ώgr`�.��B�r-�qł��J�_Y
n�pO8�lW��j�d!�Ѩ���x�'j�,8V&�`�,��Q�9�^�x�S�hi��0�? ܆�!B�:x�����9�r��,�����~����S����U8�1VRRU=�j��ԑ�C�Ns�8[�X��!B�_	��eҩdRd��h`ITM0jkf(�/7��:2Ԋ�����0<��i>7��ζiI��%z7"-d5�3,��s̾�u��F]�HAA���M!�'�҂�Ŋ �^8�ɦ8J��X���ڧ-�=?n����}�g�Ie��uU[��;�}�z�X��f���I~V��	�䠜/�CC�t#r��zz{[g.�dl�-��@^1�?��2Ό��܆�{6l޾�i����i�)Y�RD�qH��r���{&�uL0Tۣ?۾��)**����W���N-++L9�+*��R0��U;�Ʋ���4�����2C��`������װ��a/^��v�Z�4�f��(�Ӻ�3c����_x�)�t،�.Y�tٲ��O�
�w�{w2߲�#���+�t���JUe�3�!�<v�h~(�Ȏ�A���ˎ�l2�,������4�Φ�je9�G�($�ķ��L�����8�DR���,'<��i}T�A�6*�A�o��d%���'Ɠ�G
w:�3C�=����(A���`d��Ϋ�!��w���2��7�L�Қ�ǁ�޾��Y��M��luwC������Zϝy���>ں�q���������/�!z���6k񢅡`~��%K������ҕ�A�o9�"I2�H;2<dPTaq�cR��� ��.��D��/n�*�@TD�3,:-Id?�����7��ܰ�!�	�B9�X4HV����0x��"�h������x"_'��c�C�>�R��`fF����9�L \�t����o�8���,^�(�+��WĚ[� %��Ƙ�����K�:����?)V�Ig׫��*Jy%�%{��Y�f��m�
�U�y�t��P��(">0��]MM<�0�0L�f9��\\<��f4=>��?2�n��"$@cx�G)R�uw_ߴ��|q4F0�H`^��b�xPc��|�"α~��ϛ�-  �鏏�'��i *5���شk�{��ף��6�1D݈ɍ��y���� @�hi)7&������$�N�J+z���x�bL�\��:������k�l���P;���	�LoW��F�z��ﾝU7�$V�N����OwB.��;nkP�ɦ=��� 0���u&l+��a��C!&!"��K�>�%I4�n�K���m�1��_Y
P����!�`�e����]�y�~��p��Ec��"K,M�@Z|�ʥ��5��!"w^n���Ё�=��堥;�q�1Ԅ��/�'���,��4�p)�\x�B�K=7��FSW��q9$dW�u�^�`k��C��=�n��ۊ�����li��d���7�������Υ� ��?u���!F�d��s��vJY��E�TM�x��d&<8\�Tk�_m�8_Y,ۭ��`��m��`5i��𼚔-I�	�k!��\܀��H-��G"������Ao�(�i-ɢȃ/�G�eT�!��H@5�߿�|k���M^9����M�X%6w#U'���g�4����,�ig[����XT����.Qu#�- ����c�=XuO�N�t3)m�����
�|�y|��x�������w�ݻ{�ۃ|& &���Q�#c���	�$����q`)������C���B�MO�\��s}D��#,L���t�y� ��S^^
���$�v��|r�Y��S����J
���8�
�R����Ԫ�ގ�<\&Ҫ����?�� i�� Ҳ
"��&�!H�����_|	r;�l�euU��hqK��K��0[?���Y��7�%�Q��8LL����5��v�|��C�_��N5���1�B$�p2�� �D�#��r�i$� ��\nҟ�il�s�.ǚJ�&��[�t��Y�8�mׁhAQ4��#c�6�81���;*�`5�e|��ai��w��Y�/�y��������rid���`R��&zQ�&l�FC�Ђ�:��1
��R/C�)�H�,'�XeEzl؜��q��L}oh    IEND�B`�PK
      RZX�U&: &: /   images/9bab9bed-0662-4eeb-a3ad-16a556afeca0.png�PNG

   IHDR    �   �`   	pHYs  �  ��+  ��IDATx��i�e�u&��|�|�<�\,��E�MY
%YC�<$1��nq'A�8�����p ��@��#�N�@�V��<˲,Q�%���d�5�o~w>�޽����{Y$�b����O����g�}��ָ]00000000��0d�������?�%�apo�h��涿?�G�&�L��}M6n��1k��L����<*7	f"?�k�q���9χ��H)-ć��>�0�������5ٸ�a}��`1��`�뭅��?�0000000��0d����������[
C6n)�000000x�04��l�O���pߐ�B���a����������}C6>��(�!7�%o%%�l�1|X�}1000��p{%�[I�!7��J)�Ƌ�o���������J\C6n ��S�0��(�!�q`�J��ԍs_���o�ap���������aȆ�������-�!��l�&��V��\c�>�6Ð�{
��qs`���V��\c���2d����e������=C6n)�0000000��0d�����C��3����!��83� 0���fZ�>�a�}��3�C4�/�a``````���^�JC6n2� �=2L�{��4d����&�����0>0d���>��H�4΃�}4��0d���>����IJ���p��G�
C6��T��l�a`````p�q����000000�Ÿ���������S�~aȆ��������!�w=�0����������]O6�00��+7������'o��za��0D���Å{Ѐ0d�����a`p�|�?�d�N�e60000�`���Ç�l��N�}ow!�+=sTǇ�l��g������܃�	wː�{FH|`���	C6�!m``p��wĝ����70000�90d��q���>��������8��l�0���ஞg�*�e�̳��0d���v�	|#o��y�{Gfp����	#�n �C�4d��������V8,��7Ґ���5000È���!���20000x0d������{ƌ�����!���	�a`p����[
C6�sH������Ð���h�j�a``````pKaȆ�������-�M �����̹�������1�Q��a����o�;w�΂ t�H�2�d���qb����M�~fˍQ��;, �;���Ӳ�w�Bnz��9~agi�v���:�u� D송Wı�d���V\�˓b&I�PB�ժU+Oז�]t����Y"�� ��ɝ��V�>3�"���Y� �sWPO���='v-��������l���!��l������������b�9Y��xB���8��H�mg���oۣQ����f��ⱊ,�4��s��肋K;�myV�8U�('J$���e���e�e�q��>����"q,!��T�8M]������ ߰�$���t� �!��U+��4Ea�5yjY;qש�gpܖ�8��s��l͌�=�������,�4�x��&���bvv
!�!� MlK�xv-��Fz�T�U�����3*B�N��u�
�BFYEx�Т�<!\'��ʔ�WH�Q��ڙ\:���id�h�Z���_%�l�^^�I��i�V{��rQ���� ·#Ҕ?�=�y^�����T�0tp��:�i�X�Y'��?|l'�)���E��2�ϸ���R��E�v/��[� �k5r�^/M�]�T2g8��w�'O�}�i���Rq�B�5!��>��.��W_u�o���>^�����x�J�PE����:.�YO�y�p� O[��c^��������t,Q��Z�|F��]۳+«��l�N*َ�m�k��-�K���D��W-ϟ�X7�U>��<����kX|�U;���g��a�y��I���[V~+�	��V2�_�_p�VM}N\���L�.�������/���ϣ(���q�vMDi�IuU&�<��騞�"D�ٷ�@��~�e��/� ���9�"�ɥH}�7v�^H��t�������6A��Z3�f��vD}.������*O// ��j>J�����W�pά�*ȃ,-l���B칞o;vEE��+G�g��'�<O�r�D(j��w��@�"|�t�wd�,�P��d(��W��I��l6�\���d���#K�x �8*��"�s;a�{�� �G~>�J��9`����sQ!���2ŏC�V��l��H\$>v,A��� '�����cy6ND�����/q8i�8H���R�x��D��^��^?�r��E��Q���4�x�Ȍd�"�yiN��Yi��#mə��'i��8�հ�;���<D�����@��D8b������_.B��̯��m�4�G�4�<dv8E6*:����=9�3)�xo ����/����m)�`�D�`{)K�3�0�c�=l� i���%���=;�ʐ���Z'	N[^�/ہ�x�]�����H��w|<5���s�DЪK��J��F���G%�������E7���Z�o_]p\p/l���PO"���˧�n�J�lV:�ʿ������:g8�+a���=�Y��@Nx
g�H�ן�y)����A%��[�s�������ۭ���!�_:Ht�8��v����y�t�s�v\�o�M�E-g$p��[H����|Va��rs�B���' ��[��;�����K_J�52�A��׵��.>�n�&B��+l5�b�h-X��9��&�)��y����Sl[��|�O����H|G�c�xR���qm �r=�k�]m\������g£UA����o�o|�۲2|�r�V��wo�=��祸�r(
�1U���g����WI�Q��O�=E�.^Z��A�7���'�o�n�@�KtQ����o�롴;��L�M4,\A�85��^�u2[XYV���Za]zbe�<�t�q��]�p�7�����|O>��8�dW!'�C��B��B�Fq鄍���C5�𹱠���X� �m��:�_�Ϣ�.,hV+�D
R�t����a
�
�Th�>�A3�(�� ��A�c�Y�UQ�A���	�N��ؑ�R�c�

�
Y��l�
s�$x�H��ia��H�F�F�RCZ#oF��(J�F���C����א9��m>���Al�<$��}�y!{�Ae�8��t�$�y	���g8^$8�Yd�#� �%��H�C�?'e��M>r�Xd���Qw�{1$E��⵻|�4V�6�S��lt�SVt��2>�p�-�G�䁴��8t<zͲ�:|@������y���q� ے���Q���9�c�o�)� *���5屌�σ�5�3>��
_��M����#!�U�t|����� %7�����R��~i��q�װjLSZ�.�Qȃ�����8�(5�x<�<gx~��Ӂ��Լ{���ϛ��ג�kD҄�W�qh�h��M�k��K�n�<X���8��m�ux<4OHJս�sC��mC2� ؍ir`8<{��׶��n�j����aUW���]��k)���DH��8�M.�|I����NC���x͚Z����|j���>�	�Q��ƈ@��/��I�KsH�!O������%�>-�ψ���}%��e	qe�|d}�L��OQF�L�P8x�t�I%�8�����HN��M5��tl���<!��t9��(2ke^�VqZ�N1�G �&$�9�u��H��8Vgc#����l$Sa"�'#KB����g�&8h�n��Hߘ�/u:��h�}��#�KȆ�(��������;8rj�3�z���g	Ă�
*�"cŚ��L!���:@��9�PC9�lU(F '>�0��}Ty��B�ѐ�;���[=X��ak0�^�0� 5������*��  Z�	uT�@Vd����V�@A�%ɔ��*H4�<�����ʏ��
F�R�P�,�Yx��������8�~7���`���R*Dh�8!3RxJ�[����z������13@��5.���G�XHZ,��5�c�KJζHA�	��ǐ���5�Ǥ�� ����A�KhI�q2VT�~x�>yuх�����(h=����0�%Ђ��8��3io�Y9�8r�H�ɂMd�"��,���t�uz��rEQ�ͤ
�|�v&KtOlK��I'��_��Ԛ�g��ϴ�y\t_<</��*I�����HXp.h�D����8h�B+�Osg�I�������F�d�5�����=VXc�E���-2n(�|��R��sB���Ӧ>e�"K'��{��{K$��4��~jm ����eC�A���U	*�n���50�C;��?�4���$x<�R�Ƹ~h>'�q"Y�<V��:�X�d�"�� ���MV-��D��X�|}t��A0����42Y�c!����$bR��O�O�c��A�GJ��{D�����c!�ZP�����-^�t1��DNd%	�$R�s�f�AW�*YR�i���v|
e���{�kV�ܳP�9���6�77��������b����k�G�Z��/�x`�=�xC6n�C���a����8�⬖�`EQ��hY��f>9
1T�)�b�y�V����v͆������<��
d��T 
6|���&p(�r����$�F ��߅O��z�
�P����Q��R	��;�-ɒ!?@PH������%�d���g�)��c�,N~K���m���d%��dr�%e�У��D$��	I���d��g��sC?�0����Q ����6E�)F���C�EG&�� ��$B�	a�PyuH��>�؂.�2��)
����e8����8>$[Ee2%��;�Rɂ��
O���J$d���~�-���'��>��P!�Uޝ��������[�Q�^�d&#���
E��^��%����ޠ�^�n96	�']��M��~�y}q��r�{'�2���&{�y�l�
G�(���&|.y�����E%EĂ�{I�{������=��<uݴeAD���6P1�\�����ˉ٬dHU*�\2��\"_ʋFs����*$G	E����B$"9�<H(
���TV��;�9A!�c��GE#��q���+�zNπT��,^���"�Hڲ��d����ф�R�����-�'P^zn�{A�B�P�R'b(
�k�|�>ߣ���Lhc31H干q.�Q��Z��{T��n'a�OW'd�d�ɨ��<H���J�`�C$��_�A�cO�,4�$��h�X)[9�^jס����P��؀�����������ϭ��7�`�B$I2-�{��iA���U��Q
C+m�1D��F�����|���vV�pP	�(hEB)�����D�i#���N��7�sXl�0��B�ͳ��`���� -h�0J��R"_
��Y8z�18����8�\��������!x�B/�ކK�W!A˳�5⠠�Qx�(hK��-+�d�� � ȝ������k;Z@�Z����p�W
��%�à�'�i>�����-���%�d�HB�҂�ty�pd�]�)T�aaM��BND ��� ��^W�%l��G#E˒��$,�b�׳<aO���UQeJ�"a �&�:R�qN�p���PZ���D�h�B�#H�0�$����PX⼍C�dP8�1Fd��[x5��J�xn����l)�D<�e�{n`�C��s�3^y7��n��.��������L�$���͡�\rz��9!N�''`e�Qh����%H����nɊi4$��;v j������z�(rƉ7�KA�7� ��5�CIE�A9�4|NV\�O�=E��"�s��ѳ�jO�5 ,�*�.2���$�sѺeIF$8a��^����2�5�:>y���)y��U*H��T]O.ǡ���#8i.�S�-YZI+/�X9�9rs[=3��������g���u�uS�- �X:)�.������,P���
�ш�x���Hx�y�+K����ˤ���7x�=b��f*�c�l��Xy���wQ(���1�����L@��@=��<ׂC+3�4SA���Z�J���x��8� �t��C2�>��r��z1l���lL���,���sB�]&�{���ҫ�� #*�;��/�-P�׾^«��C6�"$���B��<V����E��j5�Fa���!D!V�F�:g�l3���|�k���u��&��6�T��B�0\�@�aq� ��77va�B5룠���tQYe�x� |����B^>��k밻��F�+�ՂC��D�衅�g�p�sX���c�@Q���,0�:*��ݸ)���P�tH-��K*�`4B2��5W�P'9� (������,[��b�9tD��{HȲ�(�@��|�
�	H���qn�C
��4[���ɢ�P9���%�D(�IhV��q�*MX0W�ˀ
0�k!���x_�*�:����I��sB�����j@D�s�ɓ)ϩ
�L��|��FV;���<r�.
wR��@���曔�+[�8�X�#�g�H%�@T4;	��9�zf����`��E3����)!"J6Z�������0���W�����VT��F�	I�x5��Z;x�i�������8���H ��h�d�.p]����릥E��z<w*7�,x$
*O@%��"t�c�r_2���{�t8�!"�� M�*$`+�����]}z��✔\+j"IW���Ϩ0�d�b��jG͗-&d��&ȉ��19r<K}Fd�ZS��3��| :�{�L�S~�tQ�P�%!��*"C�(}|gJ^��$��W�R�6]�*�U�p(\$'���gr��ɻ)Q���}� V�0��`6(��t :w�Q������$��Fx+��G����
<<��f����\�d�������i� �^>�8DH(LMy)�5
�H�Ӂ��w��@�1�)0d�.�����ɗ_=�Qh[1�LȪU���G�U(H�u�srxp��W_�k�68���'`ߡC��J������0?�Ċz4�n���-� -n�[h��-h�M��L6��ݻ_�.�	�N<���`��3ϟ��Q94Т��@�Ӆ���
�Q�ʍ�gA��̣��k���q9,A���U� d;��,o��`�l}�� �vU�����^�d:[YF��U8F���5WtR
2�UR%����M���P�yr$D�{,yS&l��灬1I��D
�nV`d�Q��xc���C���V\��(� �F(��E�'�����߅ 	Q�������x�g���<&^�1�83<ybK��)l�F�S �O�*Toa�۸Hu�deGă��$O�"d��g��N<��=� *RXz6�	9��R"��Ā<R���#���g4.&��l1�Jc��=��/8�A��T��&��e9�{Rυ�c���HԵ�t�����Sa�:��>�Zx���8��ӽ��C�5�N���O�9
*��$�� �����*��&,�~�"'4Ʃ��r��'���,t��.sT@ה��0ҏ��%I�P"���IȘ��������<|��h�� K��2"y�+/
y!�3��佤Dt1��uψ\�(��t�u|=�
�!{˘���j&$��ؓ�f��P6��Uh�Ԣ�!l�����x�d �a���E��L��S%�芻�j��\`�R������r8ר�+Р�n"1����J9p9��lGyK���*�[G������n��
C6�8�~�H��P�PѠE�l��~C�3p�8�N�M	5�2�7.����� ����.%�Ձ�1�.�!�`ss._�		_��)-XYޏ�6Z�dq�V_^�A�1�k1lln��k[0�|��5�G���O.��^x�
lmlA�v���	*��Se�0�F�������d"MRq����.X�{��Rm)ʝ�I��Z�KU��Nq~��X�[�0�,U(��e�S��*t��۲� /Jҡ�.)<Е"�J��PY���(����k���aPi-����`˔5I�J��,5^rœ��,kz?��ql�ymH�S؅�����1s�d�BKH�(\%r5��%M���i�h1�E6Vj�����+�n�4W$/����qR(
q׳� e��B�C_B����C��	z89T���B'o]�I�`o��
��U�`2��)�$O+k��	�0�:�
��S���w��Zt}�3F�qf�CJ�)\&Q��L�1=�@����[[� u5P�tN�gSKϒ|I'���2S��e�+-}�+I�N����E��X9^o���*iT)k�z��Y:η�q�kI�KW{*�N�7��0�~�����XJE�'E6�')������F뉼��-�jJ\��P�iA�N��uU�$��h{������I	7��j�g��Wa�Wc��@��o��R�i�/Ũʤ��s�Xk�b�K�&�Z�«6aw�Q^����h$�Q'�K��^| F���i��M�!w	�8��l	T�D� ��5*Kz��>H�l	,��b��F�砆J���0�\��\۹��5��q�ۏ��/mU�~gyu���jvQ�(�!\XZ�9n0����}��&��!�ہ�`�5�s�������q���shإ��@���"�ݭ!���@��L�"��?m*T���3��Zٍ���(��T�]��B�O���RI�R	RN�q�D:>}��6lUE��DPT��b�u��<�ʲs@U�P�,�͆�Je/G�	pj\v�j��YUf�r�8��> �:�B)&:l]
��h��ګ��?(��a++�<�T��'����z
QPf>�2e����J@�\n�BTC}�By&�b�+*��:�C!��:w8�.U�U�irTIj��(���Unu�?�9q>��n�cr�:7y�(d樔Hg�d�HUR)�^�_RvL���J�[co�T�<�$\Ɋ��Qs	�#C$�*kȻ!�r�s� 1=M))���brNFQފ�cPZ�jNJ%�G�K�\
[�&@51O<'*�8%{�軂�0�Wh��v�鰓�U���0c���h�W�8�����"�R3&.���:'��RUVnj�ӚV��$������Oń5U�J��Y@���a@�gA��F�(+l�����r2�94QԵ�4�H�(,���됻��5�-���p�	ʮG�:W���N�b��Ӄ������(�fp��}m�i֠z���kpigb+���k�M���{yAލ	����I�0d�.A`�΀JJ)�@f[^T=b�C�!�\���t�A��03ӄ}����^ۆhwZ��K�<�Շ���v#�i4����s�Zm���D��ּ�{1?���~��H��*�z��o_���m��a���
�Q�N=3�'B�wߺ�c��0���Z�C�P%�U<2P���Z-�;m%+{�;��*�}�PT1d�~�U>nVn��E�SuI')Vʃ����U�0��J��&���
N�׽
�|�ܴE(��W�n�LYRe��zB���I|�����2$�@���8����"$���*�!�ti*��S��^���E�%�P�t�K��A�%�zv����=UF$ z��"U�ꠐ�P� }?T��+k�f>�f�%�T2*Y�RR%�?��(�d9��f�o��W�3�֘l��'�,hNg$r'&����g\�W�D�Q �Ad��V�����K%ժj�\	JT�j^@-1���?գ���σ*�>�V)��^_����r�0	Q룬�p,�T�W�{�@�U)�&���%�`)2��J�\M"��M�r^�eO��3U�:lĥ�R�K�
k�>��1
��xT5��(��7ym(<��N��  BJ�+1��+��[0�����<�h�J�zz���}��Q�ՠ��p"�j��������5^r�>��C�]�3.�81�.lv��4��Ex��<�D��+py'�Ri7��2&��rr��^�50��0d�.�#�������K�ٽ˥���z}p�X$̻	��>4)��Q��sa0�v=+��Ǟ����я�x���S��T�S��Z���+��;;��N|�Vo��6��0�p���?���~�x��|fV|��!Hz.�>�#T�^-h��m����rE���^WV���.�5W*�r���ZhEYƫu�����^��(���{П�:�������Imi��v�2�ФC*�ʾM��=:��cҡ��Y@�*��Ve�B��Y-K�F���U�9
E�?b�P�U�ׄ͊!�t㿩�8i�MNy��R.qN4�%���2�_����Y��^j!�n��ϓ��@P����K�:����}X�w��
`:����B*B'K�*�A!e�L�ظ&-/�����%�F"Y��
&Z�*Sn�rT����ʒm5�S�$�;���҆��@�� ����PQ�H�uǤ��9��D�o�
Ǎד(��I�ZO�1��b�[�?��U������B��s,��PBr�	�������2��d+�Tw�d�4�匕�~����t���=O��U��?�'��-�غ4}ܿ�٧�ת�Jl�����R��$Uc���pMV�Lτ.4�fP�ͅ94�"j͓�\�%���HD���Ņ�M$��f�j��� �
�:�bo0\�{˴<��.��>�ת�_�9g��Ձ��0��U�0����%|x���[CB��~	�աX��n8A7�l�Ep��V�К衠O(�a�h�$#��~m7���=�G���e�§~��_{����~���s�Gyd�����/�=������k����'�a?
�X�~�l_{>��9x�U�z;p������j �z��e�K�
E(eU��A�p�h�D�!��-3�'J��_&��ҲS���{����D�� P�]����(�u�!��)R��R�F��8����S��N�c������K�� I�����4t%ut�Er_�+*�j�X)�x�GBYE����l�xi���<�I[�[��SI ��Z��7*Q�!��6�F=�^�E�3(&���$7����¡N����(�l����0��<��pUH[�\��s��V�@2E6TJ���ǽB4��m��O9W�i��H�l��KY�D�����Z����8K��
n"%t������V��*�27�㵀�Ly��h�!�q9��fZp��='�0�7�7��y��\%\Z�4(������"6*��+=�k����J��a�,����_��)D�Ʌ���?r��n�ۘ~ZȻ��A'�Ju�9 j)��%�B��	��5��L�9	��Q�������̈́��?54�AUkV�A�RWU<������L�cǎ�~��z������v��j�lr{�^e8��i:��u����v?����F�zݤ�։`� BYTO���� �w�wסhV�=��hs����r�����]�)sl$�e�6��C6�"���w2�-�4ǟ�������{jT�U�R�"h5f����}���_�ѯݬ1<�����o��_��z��_�ol��Yc��v
��~��?�q����a88�Bm����M�KgؕKnyU` �����`��K��/-V��\%du4�+�1c���ͅ�d�Y���/�$R��&K��<�͐,��*��8�X��5�P(�2��.=�SIv�	TwU�t�h��@aUUD�ʦN��z8o�*�q�G�/i4����-x��+\�tR�����^=��=
�;=(ތ�T�@%�`�Ղ��E� :��1�(l9����@ɋ��KY����"� �R��'��=��L�}F
�&Ia��ЂZg[�q�0�9+��$ZV�)M��H ��WO����'��G�ZQQ*J.U��e��i�Hx]� ��Q⪥�b)A2KUr+�T�փ���jMT�m���6R'��^m���
ɹ�SE�Vjin���e%[�Xя�:rr$�(B�V�^���V�:wE�� ]v.U��q�p�߶�imMex2��5�}��y�xΧ�tcR"�d�kZn����GZ*T"�ׂ[��ODS��	�"�:�'�b{P�9�*�G�=ר����H0�h8�7C��I�zl�_?r`�=���Ϯ<�#k�M�D�����{���V��A�;�=q������s(6��Q��F�V���]�������As	��[���pvk�m�N�c᮸[yL��n6ٸ�Pk��Ug�D�Y�wm�꡸f���E��z꓏��/���#��/~����W���/~�[�^�x�'� f�h�N�t�,�*MX>xVf<��nBծ"�A�Ԡٞ��݃���vT�� �N7y�9!tҡʦ�.�ڙ��t�B�,OQ�J���dSM��������[h!�+W�]vh,3�`��P�Yjo���q�����R�e�@��%��1�5�b�2C�Q9��˽9T(�=
X�p�.�7����/�����_�ӿ���t#T�u�Gay�,ǗmN:$a:7S��}���?W.]����?���wU�ݯ���ԨwD1��E+��Z�ۛWan�	�O>�}�a8|� ����2뢰��݅�x��<{Ξ��܁�0�Bd��E	�*7��mj(|RP�g�J������a�������^`C������p��&wK����eE�!�I�T���+�\�\�k�Q�}tb��J�գ���9�����B�^�j5�j�C���޸�L�9��OyG�$�a�%����k�*E�*;��*=E�A�M,��C��Vla�Z])�^�8L&��e�b�I��i���2aU/S�*�Ϋ�[��_y�T>�Nj��+wI�%Y Eʅ:�:�N�У�SI���M=�F�}��*��gu8p(+�t�d�TͰ�VC��ШV�P/�ׄ��o?�������#�؁�eq�wG�\Z_������,�~!v?��q</�59��cg��VN>1��υ�7q}��4�[�BwYC�l����M�!w�������*Hva��W�:pa�<<x�Z솿��'���_��~�+��/޺������?��/����ku�?KJe��2w=����l����*���P�*��{A��u�M{
89rl�O2��O~��}y���S�]�!�I�\�ce���*�8�͔'dϹ���<L�ī�6��ȸ�<�.3x�Y�iQ���z����i�
D�k�^��A-�P�;~^|� 4���
C���^��A:�ɝ%���0;S�����#���	��/�w_|	�3��Z�SY� �M	>��l4���Ux��������)x䑇���C'����7����^|������^~�#�̐[��Ž��%]�<�PhF�!Y�5	{�=�s�Pk6!�R� ǵ�ɽ7<'��:�Z�8�;�!���iZ�ڲ)jC�͈�њJcV�.T����+��a��&��k�u"�#*�z�s\���"j�G%�q�z7P�&���P�^U�B=\m�c�)W�d�L%TN��`�\��s�����������=kӲ�֭&b�{�X�!���wø[�[�-�j�����G���6���F����39���.̷\��A[�V��D����῅����:����\�=ǫ�<t�ӵ��HLs���Nϸ;k��o,6=��U8�T��ӻ�w����G�<6����l�E�l�<�P�k��ΈT�r��i��3�ZT�#��ɓ'��?��/X�%��'�GO�����?~��W~�ڕk�P)+�ccZ�Kˋ0�QE��.�,�Q)6��G�'Ġ�i�a�U��n�T&��0J���P�Ϊ��)��aӘm��p|L��P���L���k�mBYN���ˠΧ���*�*�J��������h7%�Q�-�D�5ꢂt`�7�o>�,Dzo�$x��yUQU ��1x8�d�7�9p�ͳ�{�*{OΜy��
5@��#F�:8�u��x������~�?�	8rd����;�a/���m.�l"1 2��O� ,�_�;�����8>
K��{#U�+��\��ph��{qe<� B�L]RG�		��x����}�<��b$��ODPs]�
}�O����^&'��<�i�d�Z�����\��n�Z-�;�v�!i���HB�U�;4��e�J	��H@���M�"R��=st�����^&R�΁I��8	�l�r�!�{0�Ug���e�N���;e�ú��7�=���w��̞�-�߄J`cnn�[r��UC�:�f��U�E�Ia�����\<|��r3��4��k��v-����������Vk��B޸�J��SڮV���x��.˯���x�n���C6�"8B�T=:iZ��έ�_��s��Β�F�O����?|�v�����<�{�����.��Q���ܿ�����Eh5]����B
	�SS�}\n�:iEY�Zz�U^O��ZeZc�?��hO;l���3>97�О�2��̿�s��sJ����W��wJU�yJETZ�{���+i|Bu���ߍ�]��?�#x�W`���C�9���Ӱ�j��|�I�EP���8;(�#��`._�F���
Zj�M��ţޗ~�G>?�s?���BIΙ3g`��=� �:�p��%XA�@�F�ȉ�?�IX߼۝�}��b)t�����ީ�7�Cet��2�.ϢBB+��v^ER0?3�CGQ؏�ǝ�pw��l�m�nm�U��6 �2iڣ�,�Ty��$4q>�pm�p��Y�?�QX]��C�p����������w���5�j`���D2�0�����Ry>Rj�li��sL螖�ϓ��2��z�b��qX�x{��=߃2Oiʋ��u[���n1}�)/"���{�3���>7tKUC7��Bly�;�ζ갰Ђ�y�Q[�vz�n���_x���� ++��^�W��'���٭Q�3y�"$EC$��?U�6��}�pl�<��6�%i���A:7�l�EhU+W��M6����>��]� �\�j�]�4�}�o<��G^��c;���������~܁]8_����+��8*��u@��Ӵ�G���,Ҋ��I�`��i�̞W�jǯ��m��K1Φ�:��1HU�@�'�����e�ypuA	j���ʤ7��f��
CN�{�+��,	�9S韶�]<E1V<<l�^PJ���.2��(�Map��H��C�Z�)ln\E��������v�ē����i����gQ�~�5�&��Ê�р�
���JFic*��������<��O|�\��O��}�����x��F���'B߇���O�>� <��qx��_?�]�§$X����أ����j��Z���/���,t�ב���(���|���Q$s3mr����6��l��~�w uBj�������n��=L�=:5�Z�����Y�va}���wa�݄�<u�x��Ά��E�;U����M$n�/�&�0L������G}F�.4�:wX���r���Ҹ���k������
o�
�%o�2���I(�m^��8/�[��sN�K�y&��+�?�Ȓ|7r���L�H�)]����d��Y�`y��J&���+\½�����?��_���oY"f��ܾz��/67�g�������W��n�Ԡ�����sK�ే��ӻ�;��-Ӵ7�l�E��гr�ny�]����|��m�EZ�^�m����8�п�c{�ѣ�_�������[�F�6�������j�W/oC���Q�#�������2,��2�`���\��uhC�N��M�ʾ ����Ke� �+]�v�9L�A�wH������({�:�b>)���x���d<�ˆ���m���2��P9&'ʒk�*x
��FTP������&[��^z�/���Ks��y������p��y��l�h��1T��B��I�u̠9�'s�μ!
�����~���7��M��?�X�؄O���#�EH���t��g����.�?�����>����$�P��L�T8(W�Th���F�����\8�&P�pl�[����U�`��)XY=�W�P$C��X�v�1���u�,���(�o�������R����0�d�����x
���ɓ�w/�:[�gN�����8,��pO����xN;@�7���D�?,m*Ge��'���fs���;�E�˝���~<p����\��C��}#QRk�ЮlV���=0=^>��x;ƥ�T-E�x�ڴ0�Dޅ�&4��M4�{z�	A���#'���%��X]mn��������|���?Skt�֨ӑ�R��� �#�\;8�޸L�؂T�t�;d�$�b��]���h�.6Po�¬��4�B߅Z�o-/,�~��w���g/_��J����桃�@<����ð�0g�l��JN�L�>�Mծ\N,,���T�L�i7�`��<K�-�u��αPAyKԾ�׈Pɖ�S\�=`��^��h7�L�(�ǒ�[1�5��8�O�w�ht�R��$��.�T�ݘLWP.	��g%\�Cg��A�^�Z�z�2Z�Mm��8�}6�/���T�M.���F8�-��;C��-����z��G�E�;�.*�7��^��^{�������8�f����3ϳ����6����0�znf�U�M���DHܙA��B�Ge=Bⲹ��1np��G4�ط2���@w�,�sT�x��Y�w����.�iF�.�]ST�,&�Q�j�M�Lz�.�D�l��=5P���5h�����܂j:煴| �g��ۆ3;�x7c�Ӯ��Kpʍ�T�T9&��\��|���*̦��x�ڽ
\��xk����X�_O��$��g�8�x=���='�F�B�m\�ǣ�)��s�_M���K�-�_ɟ��'�'����|��p�����/�����������2EK�GH�zHΗ��`��<q�\9wd"�TM5�-��C6>�D�P�Tk��D�؋sh��C�%H�9�(�g΄M����n6�9����lnl<E��hnm�s�I�ЋvN%]�6r��Z^L��#�����S�=���J���X�4Q�T��rG��7vbOJ�q�JL�un�,������=&1�h�bM�jLy5J��쏡z�3qN�.���i�M��X���UW��o�q9D�#�H��z��ų`�U��l�V���")�^m�De�A%:E�U�`��	�x�cO��ϝ�{1a��\��B��^�z�����h�D���$��$֡�l����`ie�`�ׅn��n����p��1��e��6Dq�92j�7��5��*7x:}�4o�ƻ��R�BG�̣�>
˫��o|���y�J�"��+j�	jkw"Z*W����)4[$4}�z��h+���j�a0@���=��|��}�%8s�<tP���h��� �J���0D�3�py�*�YUrm�Fq�lh�H�Wđ{EӸ/�[<����h�)�����{5ձ�qB�x4������6f���1�`Z_���Q���{lP�V"��Z}��'�}�D���Ǐ�ɩ���^x�'w�v���n7����Kbh��t���F	�(�0fo�[�{�l��U��D�3�n��������6�\N��:|䑓ѡC��A�U�����3�g�eYV!kygs.���p�"��ۤ��"���OId�^j�
R{8�qr'oYM'�R�Rh�Ƥu��C(����b��R����Km�v�z�Y	��/�R'�U:4J7�J��$?�U��X�O�4eR=L��6ZV�L�����@��G�y!9΅�Q�FHIjЬ59��-hV-�*���t��?��EX�����7l�����Z�͛�G�����|�Sp嚀k�^��z:��K�H-�ʡ������&���|#��5�����s��[	�0B�B���s\�t�+=
A��~(Ԙ�f'Ksn�� ���Mx�Yϥb}T�#8��9�P1-�΢�w��O��lCָ�ůԹ��=Xh�aj��W�x��䅺�F�!\��fO�]x�ٗ�_��o�ɏ<��/���_z�t����������ƣ�Kx��}޿��X�i5#��.���Q�?��}c�q��t�MƜ��%9���	��6bb�%������=%�y'���pɄ$o�{oHf��T>��J�^�������TB���4W���WWW��m���\�/��?z��W\f�G;0��'���9'i~6�ן67���Ð��ߖ�{������N���t�� �3��[,�f�Z����h����.����Gr���=���XU���\0�,�V\��ȸ2�X�#Ƅ��{T��w.�n4��~��)`���5i�̂v�U_@�q�+QnjUzN��8�Ŝs�vO%�Y�{���=�ބַCyf��.�T��J��H�q�[�7Ph���i{un�msc+r�?�w/���a�K��x��s�{�H���F�@G?ȍ�H�QI)]�C[�s�&���G{~��fg��[��x������Wހ��m8x� �/��ǩ�K��Ǹ��!�槑 ��o�K���}$Om��n
��A~��	�BRHz�e�������u��@�T���G`s���IP"��㥍�F���d��:�z�l��J�Q3����r9vgg�m��#yo��K�_�K��/}vv:�x��=�V���RuL��Ů@�����G&9�'p=��)(�҉Ǻ�87�e��W���4��UD�W���r��hڀ�>>��xk�����?�U6�P���y�hg]"�:���B���l�g�V�d��S�[=�X^^zqvvvk{{{����	7��Y��0���8%�Q�%����Ð��K���t���6��	n����ȶ_��9��Ѹ��K�j-���~�2�A�(���*��)��8����[���(�%�[]���XJ���$�L�Ԟ-�'�Z�=�!�f^eI߷�\RU�BCW��v�|���Zy�suŒ�}��M5��gxb/��l�5ná���I�L�Fi-�
JkJ�K�B?�h��g�"��!(�*̬�@I8w����@k{�3B+R�'�����p����Ly؃"�q��̇����y�W�d^.綬����k~���]8*���9X\9�d����6�����6�X��K�z���)ٕ�2�Ky(���ո[�7�B�=ov����bu�Շ�	�!)F�v
��s�n���P�Ig!���Z�S3����j�|wk�=6�9�]�Tg!�Rh7�����x��H\ �?��+g��� <Wy���D
��E�<~�/�w��]\������=�6���;٪���&_��,{=SLx�D��_{11)y����C����I�y��\Qk?M#(����Y8/�Dy1��|� o,X�z��ۻa8wG���Z�����ٍ�ڣ��q�}"����J�V�]���60�(� �l�%��W��Z$8}��'	Ur�ǣ>��]���~KQk7F�VK#��hr��W�*�O{U���=�-��I�H�ފ�����2|"T���E�����GQQ����e����e�%<n���w���7�*t�JI(��5��ɵ���}{��eJ�hi���Q�}>�,a�L�kG��+1�N�F�s���a{���~kpp�����8��?�B�})�j�M��*�0��1��ʛ�_zΟ?�}�e.?�0��x�o�e�E���=>��	 /Щ�_��|�k��8ý1Ҥ@n�vq��Ǥ�OT�о*�E����yh(�^��j�^����D���5h}B�1���A�����Ia��+)i�q'
�Qo��F^y����vw�^�333��w�(|�G�����ҥ|��UN	�t�� iC"&U��"wQ�ܱխ4U"q��[�C�_�����&�s5�&j0�k���c�a�tx��7�[�2�xL�x����a{��P�����0]S����ԛ�Rk���	C��"�n�R�� ��Z�r��
&�ɨ��y���'�Y�9D�&#�o̤�%X]�F����� ����R�7�ڷ�̮�J%(���F�Amn~&�Tk��wX�S/�s�'��-$K�oq��)k��`��K�1R:l���{^+�1��I1Ҹ.�	�j�('����UU6�B.B��S&�:�^�%*�Q9v�&��n���S��]$�qY���˄S{L3��z�z��4�8��{� ��N�U��*tw��՜��B��G�\�>����sً�GS}�Y��9�&��x���R�sQr�]ߎW�d����%g�\��[Hx<��Ce]eVUoVP�o���No�.\��7Q�T��]i]Pd�R^���d�C�l�ΛT��JMk��ϯ��hCF{��	}�+>�{3p��֮^T���{�� ��dV��ߤ��vF��x�PKv"+�h���Jc�b���vk��°�$/�:0�2Nj�PQ�&�ߖ�~+�=����e�*A�/W�D%þ��2�:�W�S��w�6�{ {�2�`B���~����g��M���z�2�I��N`.C����M*��r��"��	+5����i]S����M��+���W�|s���N�Cs����C�vԦ0d�t�Wd�n��Ek�KG
o��b����h$Q	ţ����:�%�u@HE>���:�;v��Y��oA�^��J�#�K�)��I_y(XB�} ʞ �-��DCy2��P
	�B�C�]e�K-HUu�d��㽤c�*�aRf;���N��p�8�ojO�=}683�z�6�{��JTi�����ۇ���o0�������3M�� �Q��8�Bkã��	ud��� ͆`�	*�k�׺�����Q�"E��A��R��-�m����4:z�Wٻ�����9�\B�P�n�J!�nq9������\8}�:�?�BI�T�5&����.���L�R�*T���!.�zP[�
Y�~�"A�n|7�=���L��;C���N._�hHyMM^�k�5=�S���PM�?�Щ��C��U�rs1Bb<���!i����9GRfU���C�
��.��^�TuC�;��s��:�^��z#_�K4�z�"#����H�����K����=��^8�[0��fn)�S�*Oȥ��b>T��f���_#��ֽn�*d��2:l��S5����co��`p�q_����h0�sV��r|@i�D�~�JJ遾v�=�G��.�eݱ-��4]Ek��djp�0�����igQ�j�2��וb���0]8�d�F�j�������nA>A�&|oS��-�&=/�-����B)�Bo���V�� u_���_/� ��Q٧T��*�e�'�MJ"bs��G�u��G�*ö�suT��*�Y�`��T������f}XGkm�\耿І+�/B5h��v-���
�0�����|�x$#9�.l!���R��M�γ6^7�no��l��
���m<?�<6���P
У]�-�Quo�dT�CF�o�d+���݁���ZZ��H��ƈ~���8�����{[�sGV:�p�3�)J�R��$�8ǣ^��;$�{�$�֮\��5��	|�J5�`g��$k���ex��������C���{Q�Hֈ$I�))0�᠁�\K��X���UvL���~鍺F����W�lG���_��L��zn\�y�[���G�Cn��I�U��9���_��yB9�9{�������,�mφ��y���Z�%��U��:D��Cj��$����l�͠j�?�?�Z��%Q����.^� �����hy6W���p��E�ƥK�*_���?q��iWJի�^kB�ц��]mU��*O�����BLż�^"m�Tp2�(� ��U�Z��0��S��R����Soj�\�WR��X�LRk쮘��P�R��A�5��+(��$��6�;�Qt/���Sn��G)̴Z���6/�c?���}~�w�l�m�� �`�І}ОA��Q0pt�����Εkp-���~���x�����{��uV���������{��bS�#���@����_~/����� �I!� �� &4�q�-˲�fK�,��4��v{=��s!lp#f�S���k������~[�-U�C��DL�c\�`T�97[@"6�T*��L%�ɥ�����`Es*�c�p��
Uj7�1�Ű[ګ,�h2mdʛ�!ɰ���-��DR�[� 5�4d'E��H*���F����x����� ֟~��sT�$���UF#	MG�e��JP���x�qW�W�k.��z�����{pll��{+���2"E$�#�5��4��k!������	a5�gM�o k-��Œ�P�)|XR����0��?��H��ʣ�a__��5,�e���i,�So������GȽkȽ#���t��2�٠�Z����\W#j��c�伣���g/����taD�~D�3*�F�F�|ē�Nn/�vl�J�ڳ�l�Z_I�Q�;8:2����x[s(W�h��=3]�=8�\>>��8Ǒ��S�g�����x��[Ka�1�/������}>�c�z���嫶(�R��Dl?$mB�|����[�k�>�#3b\0`~	"'��2����	��D�}ל[�1gk���J���;"J�=��3�p��Fh��	B��:�-���h��<�>d�NP�v .�����WʥI��� jl~��ET������������j�����lĐFR��M��h	��>�x$����x���Pc1�-?eT�6�&�&�(P��ޔ����6��4yc)Y�����h*�Q���A؏UH�R��4Š��f-�X�W�MDG�B���}��pֹO`��1d�,C�Вc��CM�[����BR]:�+����>�>��\5C�ھMN��������֗��Vġ#cz�h	8v�U}h�r�x��M1����4ʖL�y�H�s�H�Z-D��Z*A�N��f\�mmHv�VXAJ��B�O	�Eae�P�3�ޏIC�Ag$��B�Ӱ����Vx���<*��!@�\���;z�쉣��xD��+�:
sE�d�ܚB~f�tJ�_%�7k=�1l���{���Nk�[��k��Z���1kO��Ƞ����DQʗlї���I��*ٜH311;�l����E�T��;m����	M����ѣ����l���/ܶo�۱c��{����yxF���霪]��W�e�H���	H���n�#^���ŎF��
f�Ð�tCi��\�ɞ|�~��t}~�C=�J�JY�R	S7�wuL�$\�}�����,�h��{&��RP*z�xO���ԓ;Q�up��q�NJ+2���6#+2}i��,!?5�x�G�m�e�lz�i�s�� �¬�Aa,�j��_�Qo�B��b4�V�Ty$�5ųo�^��Q�h�A�rLe$����TӖ��@�#�AT��L�h
���i�����m�d4��ay�ܬ[���w�w+.�8���2�W���ײ_6�s�ί#N�I��S�d�CD+{��C�q��r	/�=���	S�Zki��ىy|�λ���c��
���I$�,�]�g�H4d<g���RhZ���@�"�+�8:1���0n+��X�r�x���J����Z�:�_\P��\�K(���"c���������Ώ+4�.re굖:�r�V. �bN�o�Q�;xx�l��N����Fc����l*H�;
n{{�<��ML�����V'��};	6^%[�+�l�>%��q�Ĉ�Z��G��ޘ�r�z�߸�w�?��o�W^�FF�����lٲ��c���>T�ffgqᥧ( :zl40��*�ru$���̱��>A|�"f���jq[�bq��B�/��F���^��Bi-|�%��7j^��Nn��`��T�a7X��5�KbcTu�4dע����}�H�e�K�����/vQ��-R��a'V�kNEM(gb��&��RX͒�Z����r�=هߘ�2e�	��91Uc-�0���#*���i�� ��#���H>o�:��@����c9$#Y�\������ia*�vUe��ݛ���\���9[UY��Jب��ƽ��I	FU�YiL�#W�H�v��˾��X�OE�ȹ��tjr��`(�\F�ç��܇V� W�tU*�Zb�"�ˑ��)�e�],�����; �D.��p�,#��#��Y�C�XnE�&
�BCdv3�`�N�/�:��/����g"9V�4�b��C�cpp�v���z�n�ںu�~��G��&��J�^�3�+�L�o�=}K����5��\�$�n�T�ǒ��Ͼ����;��Lfn�m��'�g���K���la~"�����ع���v�|��?�s۳gO�W���_;v|�l�D��&'�k\�j�ǧ053�/��ʻ�E�F�g��fP&Z�1,$ع�Hse�;^��s��� ?P@�n3���[�8�� �"p�H:�4��ȉk�F4�� E�
^�$��� \5�*g�����y%�3��K��M�s���LIJ}��O[�����5g�C��+�VE��
�ZT�uM��Z�dxA��Ǫ&���K���K��N��)-e$����刪!j�e����q���3�yr�������Bp@-��VY��B����҉�_��@����,V��K8M蟀�s|UM��%,KӔ+A�	�#�� �b����%bp�rL��Y���,�52�no�3�U儲���� _�Rc����y"'"���v��;�ӷǌ]+W�^�cE���� <V?h%�K�z	j�o���~1�I�mG����8��S�b�j�n�~�}ç�.��e�~ �-�G'o���	Fe=�V+2��<�$jn%�>���� 9r�7�+����Mk?��T�k��x��C2�߄�.�^k������}z�ӿr�����w��G�g`�;n=|�ص�Tw*�Lc._��Z��\���+���P,���D��l�n�T8�����0C�� :c���w��­�5�1�8�{BC��T^��"��EՄ�e�l��a=x=���Y�2�FV���K�\�zG�5*H%sJj�qm��zuMWe�0��%��rm1����g	���=z�Tu��İ2��jX�)�� �D<#<�%�̨Jq��V�:�)��q]9{�[l,! '-�"�����Pk��& W����G՚�a[%1��r,r8<�͈�J@��M���D :kƌӬ����D6!מ0|�jK�gl�+�D�4Y'@�c�!����%��ۖ�"�c��[��% ����y�	���`h��Y&�.E�%@%R��d
T�w`���x)��P��C����"g���w��\���;�<�q��C��a����u�1M���R��h��y��3�d�0-�-:�0Bgډ�L��V �~S�U�*���f�0�ߣ<�b~v����m���_�T𿵓�O�����z;	��kӐ��RE�c�o�J.Ʀ�ȗZ� o�^������l?4ؐAc����7Yo���,�sY4�����<.��,Y�zd��4�K�arr��?�?|�^w����y=������_�װ|�u(�J(�p�g��oz+Fg���ֳ��M�aq�����7��y��Gz�/Ҷ�A����	���x�Ͻs��
���|�Lwxv޶5]V�S�9#^�1X�TV�״�`��׊hDK�u��(��m�8���D��P����b�)5�� �\�:��\'U_+�$b��PG~��1*�n �fE���n�r|9Gۊ��(�:P	o�-"������ki8�2��T��)$m��E��(Ucl���"�聜s�^F�Q�_���<D3d#IM#D}j�4��m�CTH�"���0K$u\2�c��*r�P���x_�f�J������`����\E��\�Lՙq��HvtA:��T`{b�dq����E݄���y��ÙBQ���f�2��m���x���kXNҿ�u��8�#���"V�h$F~���Cw.�T&�*�鬌�F��ȱc������]�`�h��##GίTj�S���z�z�>�\l�s�G�e|$�|�\�~�����n?4�8	4^�m����+կ���Tw}�A\|�Y�$�}�n����y5���c�����W?7�}��;.���WD�k�Νk���{?:61uE"�%F,�#G����u�ߨ�ǿy��O����[����d?ϔ%��RnV������i	э�U{�{�*��w��%���u��sc���aV[���X��A0�牂b��~�U`�:i%�ƶj�;�PҚWW��8ջ`BK.}#�n����e�ǭ"ՕßC�&߭��.��9A?�����' P�9W����h�B�ٜ��X���c�|]y����Z�:�vp���f_�|}=�z�D����(�����!j7�bz^q��i1����u1�)��/ ���O+o��-�+�d:��?h(q�N~4G"�"JBTaE@#F�ܴU�F��'�1�c'�1�/=��G�JMD��~D6�4\��brNv=�b̴��
Ƙ<}��&�4É��~�}�N'%vH�����H�*�-��%��D���?��*�(�[�4zB)m��`�c����uXM�����ħ]6��k�����B�V�|~������}ݸq㇯���q����'��p˓�9�FbMX5\�jN;�|V�=4�ã�d怊ǲ��H�$�U��i�W��J6�V�#��G<Ճ���m���נ�t01=�LB�؀x�������o~�k�x��7o>�K_�Ɵm{j�m�\2��(W�����A�v�Y>r}sS���gX�J΁z��a���et~�x/A�>�w�m<��J�|��~I��������K���"1=>��Y��X*^�6q��aG�����x�1է �*]ɢeZ�u��z�^Q�edB�blS2�[]���:����n���g[����eD�����"��J��X-1��oSG÷S]�؄�#���Y�=�cB��;j`h�a{�D,�S�G��o�|�k�_a���W��ެ)������<	\�j�4�}}�m"��j?��*���G�Q9����c0�����T$N��2��t��t�f���0��r7X�ڨ ��\��u�qh�m��h����3=2��Ad#H�>BX��2i!)��Z�F��O?P)5�&Z�����x��1|�PZ��j�_L}���>�v�#�rbr1а�N����ZAO�47��~�ϬR������8��$�.��hR�ZU����co��L�W�����˗�"��###������slr��e˖aH�k���x�X�r����y�:>�Z�V��|�Q�7N�z�[�bל�^��huJ�=2v��#	���������6�]�xc�o�UCRӖ�Xs����������x�m�=���~��Eľ������W��G{���1lC�E����9�}�y� 7�O_�S�yD�]���X���ȁ.�4rۻ�i���MK��Pt*<~��
�s�İ�ea8�,�V��,�a.z��,�;F�c���@������ I�5<��`	Ӱ*-��%I$�i���ӲX�����\f	-B;��ŽX�SC���b_#h���P)mDU/Cu')�㦼��Uۀ'm�P�V�qgq� ˋo6�5&��,ש���n�떂�t�K�̙��u��S�7����6I���;B���J�t�:�����j����KNyv6�dT��ҀSd��(*7�%@��(�%��DQ����Hc~N<�
��^��Hfd.�e|N��{~z��y=��%c�M�8O�p]@s�ߡ�-�#���ܔg� #÷43�$j�s�6lr�"��P�j��j5�^��,�٘�\�xˏ-���P[+2����g:�r1:#��m���#�%�|}E�^�״��^�Y��	�ߎ ��-V�uϿ�R&�>�H0'��#ڱ��jj�0�Q,̨6J*yV�Z��1q��j9>93��߽zxx��׽��)G����ؖ_�wp���<Xu��ۯ<#B���0:[Ů=15[VEQ�b���Q����oѓ@�ձ5�N��tS���pci��.�ٳ��ůb�����H�1�p������3Μ��������<����ݟ|������9�9v��/>���m�����g�g���C��y�bKy�\���q}t��;��L�XV�xg�\�)MT�������zd��T��}�-?ම
�ns*�vk�B��;X�6^��^p=m��� ed�|M���B��QO,��H�U.�#q��e#?_���q$��v	i4�J�T/"�!Ǣ�z�bCK��a��9OD�J���>xa��|I��ȫ`wT�[H�p��(�߭� �z�zT�y�d�1�%"v+�)����k�)�F���T[ M,@�
9�3pP�G&' %aP�R�\�d�����NbQS*�1Q#�2Dv�伺�Z�Y��P+K?�>	&*���E^A��Ɉ�:�f A�Q���[���D��@�D�Vղ\������f�`ɹF�5�k'��R��O�\�դB�/�)2�\
�}�T��b�5{nH�n3�H��}�0�s�P?l�����PX��ZA��D��Bn���޲��M���t��
�Y	+W�]���L�H��gtxe|{�T�%N�\!��+Wr�@.��gW@Z��ݍOn�m�|�o��z��x���Kyh�o:x�C��l<��(W��O�X��4���zj�s�{`�FB�tR�E��1�lQ����ro'�(�������Jgb~$j�dAL�"h5\��ҋC���k�"����Y�\�r��7|��O~���r�?�Ώ��[x���v�=�C�?�~�������ත�.�ӽj�*��I(����Z%pյנT���{�����ΎT�dI���ϸym!m<u����2:Im>F{'��I�X��;�j�p�����Z�0�AD;�tW��b�>��x��P�^�jJ:d�7F���	��(��5����/ź�K�����b Ӹ�-�ǖm;����P/Oa��e���s����n�g�}6=�r��m�>��|D�C6�-�:/��\�=ew=�-��\��d�3G�rp9^s�-xⱧp����ۮ��W_V�{�0�s����
���eW^" �W�D�GG�m�NTĀ�=�(�d�zUt�<���⚫.U�gv��mB!_E�P�<�o�
�^}��f�f�ȣ��Mq�M�!���}�}Ւ��Ye8�~�g��T,�pʺ5X��\,[>�G߀�/�'���ˮ���_���c����NbT~�Vz�]rl��Y��y�9g���$&g
Hu-E�P�PaS$��n{p�P�*��WG�$�,0n�Y�~�jt�ܥ�������H�2ݐ>��?��|+H��(��y�ǟA6��W[��
z f��G��>4����~�|�)�5�I��iY�)���Q����=(+8t�(��(V�Y�e�W�<���������*�>���;n���Q��=�<x��O<����ڛ֝�>�T$yG��S����	�{Ɩ�br� ?=`+2��~�ٳ'���򀍓��~s��_`�F���@2ݭ����18�#v<)���,l9L��j؜9gF<��g.x|�S��������w�ꕫ>㌳��Z54?88XN��N����/;�;<<����������b��6M,Y�
��xҹ�ʤ��0*^.5n��J����az��D&���H#[Q��0�5h?mY�fU��"Oka���z�؝0￵�87�QOl��('V������3|�3]p�"L�B�	=[��A�UZI�?��S��ia�.|�?���~� ̊�<.��-HX9l��$����q�kq��_�T/�6+�_������o�s8봳�fM?��(z�𖟸������.�79�W/�O���xn�xf�a�Š:�Y\��[�+��N��
sQ��o�� �k4%�@y�k.AD��>�Y�\����⍷]mtV�-%���?w>��/�.@4)��^eC57�|>�+�ˬ*Q�/�@� >񱿕�������~�O(Q���1\{�EX.`gjtg����?�c��ط������Q��9�ZE�@q!���;�ze/����M7������>��������������
����p�W�B�ՏL_�@g�����?��Ol�?����&,��Q�ÒM�1fZ��ȥs���z�Hq�I�0O����*��h6}�,?$f�AĤG�/�(� �í����	?u��M�~0����͉ ��n�(�ՙ�V(P罨*�\�/`�S�-�^�C8�-�Id�K��HW�V�kV�B�@�!��������mW}�>���s��\s��ۦM�rG���y�������s�%K0>9�d�tWN#|	yn��y.��0�G6m��xA��a�5�Ў�y�\�+��<`�$����b��S�7R��D��+�����ZC�T��s{Gċ͂�Ӳ�V�-Y�*��&��d�d�Z��S�sӗoݶ��w<����'�R��L2���S&Q\����>�a��Z��ڨ��[O�z���[]�V���N1���������w݃�۞E&է��B�y� p�KR�"f�ͦ_
�a���ܾ_��"2܂�,�` /M
�!�2��e�-�}�~5�B�;����10.�z�^�}��(IU^����{;n��<��|�����ø����g�P���~������K�oU'�ZqL��<�,��L5��܇O}�s�_և�����}��8vh[7������w���5��U,FP-�ѝ�ᜳV�u�P*��o����rlۺw���b��p�7���Q�{~��韼݊�7<��r]q��)�|`�%!��������`����}#G���[ߊx�Aop��g�g��6�j��ů��6�̳Γa�R��;׃L:�����s�K���DQ�˽Mz�����f�/}Q��7��\s奘�)k�ɼi���Y�r]o���-���{VΓڠ%,�r�姢����,����	�q��E����Z	�����h:�D�i�����ǯ;�J�O�PKn=�t���mB����a�$�I�'��[���L� rю��XȑR���+���a�P6z2^�����+U �o�"�'Dp�)�􌳕�[���͓�3�[�ȗ�r}�q�I ڵ�����]����`����Y�z�^���?���GJ-<���1��5�����=h�kv����b�mͦ3@ FWًgzvS����SN�y]��B=�$��w��V�/����T".㬅j�do�Wb;�Fy�l��ךn��|�D��?jлb�+_<�##(�Ϣ�?- ��<��^18$pV��U:�бF@G������[m�)W����1��DR�AV��\I��tK��@��G������)p�E���/O��7�y7^�{@'��@�X<�H�HʲB�-H �BY��b�j<�u�XH��E
߇��_7���#��au�ݎ��c[\zh/ �-�Eo�������q�^@��M5�mw� �����k�Z�`��^�ab�(��ӟ��;wɢ-^��_A����.`��lx�Ͼc������'�'Ƒ=HR8�'&���aTv=��%	����!�|ۭػ�jQ��߁}�v��.��G�=�j�r\p޹��.t���wގ^����?š�G�+��pL�.�8k-n��&���?�3��Hf�q��*�^*4���Ӭɍh�HK~?�����/�{�>s̡
�����w0�;�����M�OVp��w�'��T���54O��_�i��Y�b)�<g=�l݀������I<���Ri9G�C��ç?��;r[�ڌ?���?��~/&'�O�8�ԕ��u+��z���搑����8�r��[@QG��G\@�G���f��BV�<KF X�n�G��/��@?(��I����SM�}^����`ܚ�#{o@�I��ຣ�Zͩ0rb�ѺA(%�b�tG���K�!�
0�vr6�K"?Y2�4�l�Wj�u��-jý��^��ຓM�<����y��c#����NΏ-Y2xx����w������'z<��T�����.��.8���rϳ�d�gyrU�J��Z�sŒ6�\��T4_��=xb�Ө9QՐ��"Zb���d�@I�����������ͳ�q�ސ�U�-.Ҕ}�
��PVYlf:;�/!��K:�$
�&Sy���,��a`�u�;- ��D4���!7�⌞��S���{�`�]�����;:r �=��t.��J�]s�<;��7>���)YȻ�s�`Z*_M##ڙRV@8b�m{���.\�(m��͗.E]<�����N���9V��;g�
�X�[��1�f���`�;�c!��Bб$��0:CӞ1fw�����R����+Wb�%��������czK�t�!���?��k��-�ߊ�����x�Q�LU�<EM�r@�i�o؉��o_p����N���uǓ���~�y�l߃��O��ek�{�F\�e+W�/|�F�ѻ�T�"��T�����	�C����|V����V��&����cQ��d�R����ٹ���j����""�1%���כ��g��֝O��-�#�Ճe=�P,6�:�".���JӘ/��m^1�	#���r.֞�W_{��G�̮��<�B�ncrjZKv��<���㚫oB�@��:�^-n��zCo_�]u񛰪Y,�㷴���,�5��
�J�r�$�&"��X���(9JSĔ��Km�(����c�d�DBұD�|�����Y~��D� �g���y�
�d�O��t�h�-� �u�^P!�0��Jˤ�`"�]b�j?$��EP�H����Zh����Ocݚ�:'8���DJ���e�`��9�[,�177/k����Ձ�!���)�cz�Vo����󚝟a��b.;�\������4�ܱu'��U�\;�P��"ϮU��vI�m�On/�vl�J�f��W��"0����Q-+"c9!+Z�8��Ӎ�P�Eף�aV>�A�B	缀��j��N���4��G�5Q.e�g5-P���口\��ċଳ�G�LZ+�o�~�@�T�}�Q�R�:��R\�mzp���&G�Y�J:�&/����
�&��U�+����^�,7���;A-9�r��b�zj���	[[��/V�w`2�~PJ�����4�ƙ4���>�xwF9�/��h6��a\��{g�y*��)��[.$���.Û��zՐHL�����>�\*����mx�߈ٙ�*k��/��&doϠx�c8�o?n����Ic߁#Z*{p�0z�zq��k��9���˵Jd˖�X�zP���;�j~ۅ�d��i,[�LP�XT]�;����ē�V�������<�`��gv��w��[���_�g�}�w��9.��A5S3�y��US�2�MS@�I�Ÿ�����Ћ���Bib��>���o��/���p���¦O���fgg����'���l+_�kbl}}=b��a��\xޙr?�����#���z�{��X�`��z��ϓ)��#qO۩7Y��3}�9(���-��TE�Zuql�`j���&�e���@:�Smb�aU�ʸ�&�ᛜD{\[A%���1߲��H8J;���Ģ	�꛱�%��f��Od��~;Ja�I���_W#X>9+�g��5S<��4=W�
ǒ�6��We�׈���$2i3�3����3Y�Aq���K�/V�jU�^W2����+L�h9.�x,��oXb�������r|Y�ıZ�|9֮?{[�ƆM� �\3��N�\w쓘L�溬mQ��jԺqr{ٷ�`�U����[�6�l�HF"װ���9��-6Ӓ%�K��+��P��´x�B������L�
������.�<U�c���`H$52ѓØ��45<+^��}e���i��I��\,s��TN����r>4Z\$��!��X�H7^�2.���4�`�j����et
B��bhӲp�M����3f��7�1�DL搡�r�4��n�B�.�q��t��f,P�tL�i!�q��R��SmBA+K�дLS1+l�[Ę��b���px�Z:.�`�*ߝJٲ�v�s�i�D�,���^��N[!ǫ�vd�0< ���&�����{�����L�ܕM�Pl�R�P�g?7?�bX��n�Dx~�Al|h.�x=nz�8���0;7��c�q�Wk:!.���$��ݳZ�Ș�xd�,+V��ӹ"�ΒA._��뵦Fn�z��w���?��\���;o��w~���m19�ك���ZkCC����V��%.���:��޲0?W�1�Q)�����Y�t㕸���q�o|������G�hNc��@܇',Ǐ�X�c��u��UK��p��a� ��_�ܳaۼi׀f;T�Lƻ�p�DңJkS���kΫ� .�K<�rMnwC�T<
��m �bf��V�(�Rc%f�nS9W�"�>Ѷ\8~� �Za��y������J�DлV0v��[�.����Y�j���Q9�-����e���|��
�z}|�=i��R��4�QO&��$5�?7�"_�������3(̕�ۗ��D6�AW&+k�%`�u����9��H[&g��Y�X��
�"�nCk���\L���7��ݻ1" 3���8M*T^A�dT	׉x�J��D�Ҩ�qr{ٷ�`�U����4�N�J����Q� 	�^�ӆS,�d�-�h-�ղQ��Px�F��\� �������e1,F�\�~��F���Ǌ�p�� �RU�C���Ev��14��G2�I�L��#�$"1Ӥ��L����a���՞��M�+'� ��v��86��V�L�ɱc$�:(�6���ٓnA��H��қtC� �G"��]H�E���J�f�U�SL�'�����1��D�Pa���Ц�3#V����v�l�l+d��#�Zq�g�r�>�ssb|��+���B�Q��o�� ^����/��K�C��BN�����>����~�~֯�����:����(���byj��F����� ��.��sظq>��?�����b�Z|�o��L&H��X60��\���R����s=>�ޞ��1Kr���A1*r?TsC��FV'$��kj
�!�����q�@*��������3J��Wjȥz�����q14blݙ���h�Q� �b�N��LW�J�w#�nو�/=������o�
��r�x�1���唋��Y�\�R�P.���H�S֡���� �~(D.��b[XlԴb�vY����Y����V�;s�1p��O�p�����7?b��4��S��.�f	h:�^�Iי^$V��;�,�u5� �����vu�(�����S�_� ��n��e��f��[���oX:�MD1�~�W�,�|<��lv�^.����0�V4Ƒ`�ll��5������i�Ѵ�Ǐ�疮X����T~�����U��`p�R4e���x����e��8`2������/��~�k�[�������:/������$�x�l�x�a�1��Z1Y>n�gL��v���Փv��Qo^�/��)8`�����ˉ��	ܔ���;�1����x�F�=��a���yY��L rP��QRZI�V���1�T�d�#"��&��hW/�$�xxAd��o����Z�G�������tiº���/���m���j�J�~��I�6��G�|���pMT#�� �~���<�Jq[���z�nG�]�����aԁ�w�x����>ҋ��Me�Ԗ�ؿ�0^{��_����)P.r����O�͖v-���p�p�՗�ꭺ���M�8��e�cjr]~�>�l��(���&�I��6��ܡj��\~	��'�B��ġ�#��-㬳Α�}G�Ҟ-}�9t�c�s�U%��/��'�A~v5n11lK�(V��V��;4�,��r}V�Y��q<�yn��fgq<��6��7����Ė�ۑ,�K�� ^�l���t�TB�2+�#㹬�,��riIy�)��By߽�A�_*~��>�˯�
��}��k�xZ*ϫ��n�Z����ȑ#8���0ԿT��F��ʹN����3��`o/*2w�&	�&M���(OI���5F�l�`�$�)�;4L7�=}��Ӊ�|����{�p�hI��t��	�a*�
�1��:ߵr)Br��'Y���/�O��p3�e;�����-Xc�.�q�R[�w
�d�5��Q;��4�Ir�|�v�D+^����of���j���ٺ��aJ�R-�\+���˖.GO_�<�"�2��v~>�B���R�*����9a*��^��0���z}��PմVu��4r�7�@�n��߃v~r�a��`�U��Y�:�9ڹ��1��4���!�k�㡋��7��2��M4������L��aG%�􎠧������M���0p,)�T���N%h�f:iFtM#(p�ۧ�ELkv5���jhP�	4�a�_'xQ��9�zvV��)ILs���0Zb�����E9rn����O=�0��.��������g�s.L�P�,젩gEF�af�Y���iZE��S�⚨s@&w��}� Bz����V!��?Iϯ�wcc���羀���_�>�~�����u፷���?�sX�dP�QZ G�xs��/~�^vrb�<�.<G�S���9�\�������6�4d�Mf��w��ز+V�����p����S�7���v��k����<��4u���řg�æ'#=�7��<��y<�k��n\{�Z��C�p��Q孆x�K�3?�nk��A<��w�[�
�_y�J���Wp�}�򫯕k��P�_��k����v9�4��TJytw���_�{Y���n�ۿV�]���c��+F'�����84|$�w�*`�F���*\t�طo��g���G#\����;߹G���]��{�����a�fh��ȤZ~K#u�>Y2�8/�����B�SǤ*4�����R����VZ�����L?�|"�A�c�ʲ�ԉ���xP����3�S)�[�	:��}�`%TU���mN����0⿈�a���#�6d�)��(��QB=��lfh�'\؀�4�3�ʤ<���ϗ�7P��DO%177�Z���bז8V�D],�	�m�P(""�ee�J��
���?��j��Ѹ��#7�k�X,���/�pr{Y��`�U�Ʉ�,�Uq�~����Z��F����g�~���܀���РYL�#b�I�>�ZI=(5�Ln��DЙ��Ё��F6l]�A1����I�R���ad�4�Rނ!��@FS&�p4�˨ED#�V8����7 ��LD���θnӠ���0Ho�xkt�6u�VA	T����UN���iZ�0ϋ�X��	k+����y&{-�,����r�
���N�^HX�!j��
F��ȋqA/��� �cZV́��g�s����R�hɳ`i�͏������&��x�uS.�c�.|K�O���u�%�����eq�%c�)���׿��n@*P(�ԯ2Wģ���n{�x��ct|ٮ;:����?�k9>����ͷ�^C�]|>&&G�������-����?��?�c>���u�`��=x��徖�?��Y�M�Xk�}?�n�a�gٲ%x�G�c�3���ė�����w⎿�#�?tg�z�|f� ��q��~�G7�C�9��N���i�?���o�>)W\y1֮Y�/=K��M7�$@��xr+����+��>��E�8��4���{�E�P r��`��-R5�۶���I�Z6G��T�[K7�� kZ�5�#�V�-�rZ�rH�5(�7��h�Σ�c� ێ,Ф	ˬO�f
	�Z�����[�;#w���D���G:Q�Φ�j�F��)1;Kɞ���ʌ���T� ����G��!��Q֐0j�'L�d��q�7\[���ʚT)Ocr��}/���l�!x߹1�:vP	��Ѩ�*�
�Ҝ��M����D���6��)��k���-u x��I��+����F�����L�&�'#Lh�!F���<!'J����XC��w�pc��h���1�N$��#�ϋ��ʁ�F
(/M�^E4jZP��e;p�D�@����p!�ik5��.>�TZ����ד�N13��:�߈���?%bjS2G�bLQ0?o�0R�����Pw ���L�a��nSA �I�wؾܸalo������+~��ɶ�~Ы���"�2��f�a�C�A�~X�h)ٕ][[A�_!���jit�cE�4���z�ݵή�Z�C�����4�>���%���o�.�j�
��Ɓ�,����V&���S	�Ͽ��<�Q@��~O=�w~cߴ�3��^!`$�r���t�\/�ܲ����a�1�u,[���;��~����7\�3�8=�]��?}�>�ccc���я~��r�:�,���];�s�3�{����Di�ɿ�ȑ8����+��(v�x�RU���%���u��4x� ��y<��Ftueq��gi�ɲ%���h�ͳ{��P����ķ����w��k����<&�{�G�~��7��o�[�z�v#޵k��ʿ���g��3��ơ��re�oPK�G�c˓O�xp��n�bEEK9C�F�����G�{��I��<�/�-a��H&f$�`J��c�N����
v�rW�3�\�V�����
���J�oR{j�a�<���K�\k$9<C] p紜6H!9�
���k@7#8ZQF�nk>��<�<	*��xmӰ��T����S��I�*�ێ�W��F2MT$L��r_�'GӘr?�5G�.n�LF@�e*���8	�v-��Yl�����2��Z0��>O��H���h9n�|�愍���H����6��?֗�(W�9��U�KD�@dz�G�(±[�^aC��PA�*jsy��;��.q��h��H�32wlm;^��g�c�9:�Yab��o4͗��Dh$ii��'�pi5�e�=#e�{�� ��R�H�NB�y>�� HP��stA	AzD�oB�<oF=B��4�8�*"��v�5DӘ��R���ҩ �ӕg�^",���"�4^K�ZӀ���{���)��8#���04K��N/ˤl��E=K�0\8�@M�������O�VS�9��`n|R���UZ��ƅ����������x�4�\3���رQ�zz�^���(��ֲ��S�����۱}ch�NS��F&����b��r���l!�u�&l������11�Ө���X�J����[��f-�q�l>Cӽ}}j��2��<zd,?��w *�en��K-�H��n�{�(fq�}��Ǹ7�C�D�#������4R�(T�@��gJ���"�s�c��s�`�e*j�H��,��-�|z~�������=r�(&0Q��O~�JT��*W�
l[�������k��E(�G�jx���D��'���-��-K���K�-hS7F��/:Q�?������F�T	H�I:Ȣ�����TK�V�&t��C� 3=N�v���ڜF9_x,G#p-'���Hp���y-1Q
#��Q�&��h�`Iѷ�r��!��-Fh5�d+��h��M�zJ����9���4��-�XJ�Wq�4 ��HoC�;�y<A��\cX�M>��x�^��$N�Nk����m?v�qr6ߍ�~#�*����)��k��� ���;Ӆ�,f�U3�����E��,S �יzqLUB]���Ç�r�2�]{j�r�R��B`�.�5��Tz�+���Ѽ(��3�kZ�O#��Ӡ��LȢ�ź\�hX2��ʂ�����E-�`�͸V*Ԫ̽ב�ĕTʅ��i��M	���kNW�7l]�J't��j,�H�)���N���u�ڨMB,�O��ԅ�a��45$��ih٢�9G�r#K������ڰI#/ue�[1���F{���kyA5)��mL����ߙ����I��L�e��"�6��ň����+����������XD�C���xZ�jt��X��F�O��<��r�X�D2A&�1S��4��b>�$_�o�=��:�)����N�H��3���BqNK��b���Y���ا1!�1Q6��.BQΡT�q!�5M��&Ӂ�� ��ʓs���$���d\�e����|+�"*��N������ͪ���M��=O
��1�xʱt�XG��+i#Ar
����O5�tvJS�#G+�f��V��UJJ�ds��T���㨥�=t�i�ZM���O���e4Ry#Z��5�(�>}�>�� &z��a$H�ލ����Xw����F���%CG�^���F�6eӭ&��<�؆K�lO�Z=s���Ȃ�N����ʼ�����\1Ϥ���&K�m'<� Mi��ḌFTQ-�#�L(�`�?^�Fgel���n�"k*�Jq}]��I&�]$@C�J-[1��2Z+���"aS�4���ت�8��/찉O���q;	6^%[�Y�Z�c�^���k�5,�di��!����ǔB�\
CCKT)4����oF�OR&e_o���e�1�
��~@K�n�����L2ы(-_ߣ�(
�����'�T,�MY$�5Q���l�aHs5�7�R�Q(�&^4S<YF�\Z��k����DT
��'�N*fr�7U04����=�/_���R���;�)���.n��� ��"��K����x8��ܟ���e)
�h�Rҫ)��5��h	���"�2ylc\����-0ǿy�v���Ú5k�(r!�����P#��ş�ׯE)_��ݻu�k֮²�����9<���6j[����x�%M�%�6�{�*���þ}����{����I�G��$Е����<�Ҍ.��֮P�,�\�"�`��lN�Y@f#j�:�82���� ȣƁ���9�-���=���R��*^u9h��K���"	�<��F��qӰ��(�p;�����bPd<���
`q��U�E��MjPX��wjw	60�y�L�@R�{�IP�k��'�Đ{���Z,��8�!Օ��Zƺ�6]�
ēq���,�3j1�h��n�:��J�F:FO<�n\�`Z4��R=�WpO �j����%S8ƃ˺-�P�q>�e 'H��T�s��9���.}��&��k;� jh�%$�s�3�y�()��e@�-S&�5b1�^�������� I�(�f	u\�(��4�!�;t$lM6�\x,r1�k���:�P#EK�=K{EQ��:L%j�LWY#/7;e�/��J�ZJ����-��\&e<��r�FƓ��>�u�MO��=�N�Nn/��* ��Y/�f�7��G\�"��.\'�"��#���������Ǝ��}ϋ�PEW6�'{�0�O����K��!z��q1<��pS�<���qzj^�8��B���͚�855X�g��Rb�ȁ�eѤ'z��/e���k��Y�E�pfT����RQ}c�)�^o5Q����ggMǈ^��U������h�F�^_S����v1l�k)��������&s
�F����RK�EG<L�t.��#+鄹�\�y������� ��t���'4�����j��?ITkT��ό�W\��h����Q�&�|�Zm�y����"���P���eU<�����g�{�����G��U�$��Y��Ԫ�fZ�4
e�U0z�"L��i�-$S��K#E!/z���k1�� 5���ܨ�Ԋ����Q�䣷�0�T'�B�Q�i���Uѓ�Y��ի͘F��("vBNLs�L�m5� �bɴ�yD�>ed�+���k����-F_��0#�'�h����d���H[��Dc���F�^ɽ���ku)=}��Z�hK�@b�E�:h��3�2*�����9�Ù����˘I�!e���gesq�6�5�)�1�hZX��
:�{p��vu��q^�s<��x�	29���&�2��!uH�AϾ$@�"�<!瑐s�˹�d-��|���[����jI�uW����B�ڮ"c$�QȖK礮�^U��>3MƱ��͛�<�s�g��T0Íj�F�N i�j���Z��嫥��Z51`��ri���Z]]��z�V��r6X3O;�t�O]��܄�?2�2�ק#���J��Nn/��* '����Ly��%͝ψQo5��:E�zf;�p��qᅧcbt�����a�b1'^_=�Y�l���bl8!k2��e"�
e���b�,�i.�4�aD�;ׅz��='R~n^��]�����X���4��Q�,���e��9�^s��� <?ӆ����C���ȃ�Hh22"�L9QА1S�LZ$���n�e�>Id�'�777g*3���H{�	�h����X&|n)A����\[�v�:�51/!#���[�����ɄU��Вsqq�|��<�劦���rU���7�xN����߲$V��eňxڈ���>&'�Uj>�R�I�M�%��_S�F��1b��y(To�^�J�x��;�'�զ8�C��4�9�s��"�� 0*Ɵ[m�(�Z�k/ꍪ>7�6j�Dԟ�w�L�Z�i �x�$JF�O�Nâ��n"J<�*��GPa#�0��FĈk���\9�4��KTs��
Lro$�|2�KQ-g(���F��3F+j4b�3^t+�!���2,�B,��rQ[�s�A�=K�ѢmB�x�Y�;�*�EF��^����j���!�/��"�-���|�xe�Oϋ���X��[qp��^��3���f���	��}�8�S��`[��-�T@Ê7�N�ɸ���-��iZ������Q��)A�R?�i��z� ���wF�����Z�ajȎ�%� k�
�m��X�Ê5M�����y��k�����F9HT��U��Bw�:�4�+�{��S1�?�}�_��*���阸�˱|�)xb�>������{d�'WF����I��sn*�6�p�*^䠇SOmZ�u�x�;�W�8�qKGb�e�>KB�g�fb��7v|Gcb�؏�Y1�-e�W�48U��E�a8\di��
:<<��Mڃ�M��pa!���I�����P�#k���� źN۫
s�\̸H�Jyp�*dͥ3j$�~S���;*�ş��P�-O�/�{!�F��j�"�ͤt̹�s$Z6P�EHY�<GYd(���'ԃK�ihIbU1+:GKS��&1!\�j
x-��/��%��xY�m�92�����,��z�ʅ�����U�N~�U�x�y7S*lcn&otNbTK%�A1��J�ɨ��E]�[UG��$vzQG�KC�c]�a��GU��1eŮ9��5r#�o�XsI���v����T��j*�ƚ��|���G�`��W��%��M��MU&!t)tsMΞ3v*Z�@,o>��L<V�~ګ��K��.�V�c-mH�ZE����3�>,Uy�S����B#7�4�߰�p̌c��qv;�@104�j
��� %6�mi~�A�`;h,�h ^U�& �-V�?�-y��bp���&�A�F0o��!���oWU-�=��FP���Ԭ^a8�2����{T�6M��X>>:�.�6�5i��|=3i���=�r1(ets\m�f��bA	{S���2��,n~���t����f�P�h�3r�?�?mt2亹?'п�&w����Ñ���xF����Q/U�y˗�V��=�jDT�nl>�:�>m9���������֒����|kӟ��[�;V:������#ܻڊٞ�Jӊ�Z���>���H6K&	��kQv���5q�b��.V�0�E��e[͈�⚱ֳQ��H>�2ݓ��x�,��G|�N;���ȍLD�z�r��o��x��X�7�=������`�U��i�n��c�f�j�cvp=�>=<������C�Θ2M�X-�������ŀ�m�k���\l���qS��zŔ�j�\D�]Es���*?�,t�8��(֌���-��9h4X��|��|"=�f���	���u�4�{�_�b�[T
U���R�,(��VnVLy���B1o��c��B�Fs4����0U5n�J]L}��P�.Ƙ���@(+������M�I�=�n�z���Po���F8:��8;��y6���cτz�� �������zS�HY�/�&�ŗ��VbQJ=�H�$�y�^k�jp:�O<5KT�;�<��VQ�4i,�V� ��C6�#,P�Tz]5a}���@Ԥ��H���AC��iw�=b��[(@i?7? F˔���k�}�5Oˬ	.U�Ru,Fe"-%���%�V�&�
���7�v�F�މ��M���~KB�)�v���IkiiK#3*d�]������eY�����-�&H�)H4"+�Ѡiw.6)����hL�2qh�ՈӘ��si�X��a��M� �p���F�⩘FU�L�����%4c�����������AD�����U5܄~O�M��rn8g5�'u'�q%u�A7�7�3JL�Mu���S,)D����7�,h��y��7���N卥��)i�U֌�Š��jݰ�_\��\��*�.����D�&v�t/V�X����p|��v�ͦl<�H�֯E�)�'Brf=��M�>2�Е��y]B�1U|�,#�AB�su����	�%�M��p�ko0�-F{-fu�[r��%aǵsn�c�5J1 �"�8�Ǫ2���&�lz|�w|{ɺS�Ѻ��������͊:���7�%��Î�w|SN�U�R�[�K%Q@K�@P�Zi��������R��6��A���]sf��|Ýb����;���f�ý/^f���"���&��3n�yZ^��|A����\�^�=�O^~�7�A�JR�d�5�H �ҚO��v��A\�N��J֮&W��
��"��u�H�8T6Yg�쬈O\�O3���܇ZB[/��B�`M!PZd�,k��l	n8k^`����A�u��A^�D��	��S�,m<�9/��Ţ�
�ۚ�<��,uՀeNbt:%6
�J)�}�|��}E�d��Y����ek���*��q���X4��s�	de�?�I�F��5rV�bk�e���t�$��(�=��o���e�9S�ɏʗ�մI�p�����_�y,�9���'��"7�q͋�i9�ˢ�a�|��$���� f)Cx�uUQ�2�(�u�	��٣&qu�ډ�^"��>��;�g��\J0⟔�b���&EJ�Ī:�͈�u<�p<�F�ԓ��V)�|�f�;㒐�$"�P��F����{I �h�-r��9TX�N�(&�".>��c+��6�-������O��Q�l�N�	Y�q ��̬qf���rʋD�5k%�}Ɍ����ʀ-�Wd�ź)
�Cq��ui��Y���W)���8� �c��G���b.EF�M�w��N�d�2j(R8�`TL|M��$]7��e&��s�؈rÇ��;3^JQ� ���BzE��M~��%���_�ۿ����-�]���vS�/_���M9/�9�Z67JIף2�u2�Qt7)���Q����X$�����Y"���z���2l�!�}�+����(��W��V7u]5k����ˇ�_����������V����-v��j'�q$����5]�,�o���,36���7`cS�5!!�)��r�$I'�dN�t��g���U�զ$xb�|S`$<���b�3k���ɫ�E�Fyiʜ�+�SM/k���Y��� \�7���	"~
�4��a�'�@�ٝ,�`���+�؉�\J�?4fa%�/E�e� �xL�*���7|�>�@r���S�	�97�͈ �n���$97�
ة����
��7���E����eT�h�=;��Tӻ�P_��C(؇x����T&qP��B�z�Y7�r5��Vٚ�,�tWߒA�^��$�T֬g�,�����+.�
O��Ä�p[�)�-�>���GɑV9�QU�q�ΧSr��	�C�s��ٟH¦�*3�d�|���zE.�P���X6�	�w0p,�2�ށ-/2��Ќ
�Λ~E�t��z�4?0�	nf�<�}�V!�6\���.�l�P�)]�x��6r��ں���+AeZ��*�;A>^P��\�gs�% ��{� ��l�f�
�N~"��NrDĹAQ���_0�碆�K(�=<(�(���[�³���pR1�`��(��28�b$� �I����G�h9[Y�S�����n�ke��f3e�]$L}���'B�|�07�D�������8:�цJ�r~�Y�.	��U(NE�4�2��`�XN�O���>�t}/��	<��������A���'4�/�J��\*��b�=���.�(�CP���5�%@��,�ib�Ǌ��<o�`.�Vʘ<sxO�b�S1�hѬ;7s������������ٿT�	<HV��6��*��NJ^�	��H�"���۷$p<m���}5,�	�eٴ�P��̊Qp!��H8:Q����wƚ�jbپ�~����H�u"p�ē��#p�E�:��h6��7b>*�>��+Ԓ�yֺ��M�٥����m�TocL�J��)�����0����P�M��2�.�2��Q�&�E@IU��`[V�nڈ�k��i��Iju,hE�;�E6`�������a��������@nZ� 3����Ɓq@�dѼk�_�!�sY��ų!7��f�+V\mPc 99#�N���Hw�d�P��T���ތ�T�\�~��1"�h��1�T�����b�;9BmLR)_e6Ǆ�cJ:%��#[��&`T�|`���%G��q^R�74CE cO�5�]r������ci����&�C��&�m%�`�'o]�q��#h�qLH!�# �x�gn�?���،����Bn�E'Bq?2=�w���!AQ� 0�j_y��e�"6�`z,�TF�z>٣����26]���1��B,*i3׳�_$k	��C'ʈY$R��_��IieM����%�S�27�ks��,'�/9�`��	�G��%麡�9�3ҼRlo�
�Ͽ#�6/Fk�3T<n�s��[ȯ�H����CLP�9~L�9e�/�%|X(��U�.�*�u��P_%�$�F�dE�9�	��2����67t��@�gS�jY�
�ݿ{�$x��Ƒ��*���Z\4�z�,���yM�9�Y ��ȳ7�}[�J�O'�ϊ��s@IR0�k&h)�a,���٫�e�ΫYDID��O��ך]~�\"���$�%�u�H�F٬䌹"B�J�Eٳ�PY��;o>ǃ�)�7%ㅬ���ղ��7���[W�Rb�6	/���¬�i�I�D�W - �㠨@<=�&C�ɡ��j(ʥq�ف����pC�z3<)y?]���T)�(��M�+��p�PYs�+�,��"�f㥷g"��q!���2�+�cC�?kz��)s� ��jy�@X����6QI��'�)?��/3G��� �N�J�[��xceA ��� �0`P��G�TUq�0��H\��)��1�����@���"��8�B�Ƚ��yL�ׁLF��-b�+sW�R�sp�o�e�f��822�+����s��9�c������K���Ty��qǢR�ԕ	AO�7B�����&|<nd2oL`Fi?����+����)n�6N�R�iXn�_�B�qc�$K�N��X.����1ϳN�,0��"� �Nⶀ"�h�G�X�[�7���

	��9;�`�|�F���Ü\
�-�k��
���(����~��s�075Y�o��"Af"�������d<��9����b?b��E��5E5@(CKh�X'g�p�}^"������7Ck�������6N�%]]����Z�ƋE;������7͸��H�
$�f}:Q�
�e�;�ZJ]6(�u,%�X��<A�M��J����Rrr1�]u9�ݺ���1����Ƥn����'�U{b��x�V��=���#��"�h�U��B�3D���q�~�-���@�*Mt�h�8nF�+�{n\�������Gt��\�� ̄.���N;�R��p��D%���� ��%U�H�Uw��0�~0���#3�%��⼋�� �.�\�v,���Bx�;A�
~�>k�ygCU��%��E8tbVK����"}�Қ���Υ�5H�6w��5� �{q·ʟ'���6xsƺM7��o���w�_K$��D��w<�|�~�ΐ3�d��@-��H����
���ه��!���e|��%Ɋtw�͊b-��1��Y��zFU��Y����f�`�JS���|���lƀp;R�B�9���������G���QlK��b��r	��Ƒ�Us�͓���;l�X�ւC��$[���a��M���{�w'.G;�Mf���m.�{bi7�v1�3�S�����+��U.t�k9Us�ݓod�r6�P�X��Iyʞ�Ţ�j�sM��Z��ȗN����=�aXN�i�vr���z�u%�����[w�@���n7�8��N��^�7S��Xӝ�pt/��[\���e��U��#��ڀ�6��zN�S�/12~s���ݾkA(���.o��&�o�S��Āf#΁�� +��E�	ם�Ptm_�pd������l��eQ*1]���/�����vJ^!n����?��ܙ(���cd9���;��� �e�T���45\H�]�X���Q�%.:黼0�E�q����Ҭ���dm���Q9��&�xPfQJ���"��5���v��K�A,m;����MyԢ2�u��I̻ �,V�߬����6N�%U��%����3Ů]�8Q�pfl�QY��I?�ք,��)@�,��t��Š[���p8bdY���C��H]Dl�-�^]beJ;Z`�.���.� ��#��&`[�������A9ki�_�';{O�����<�\l,��6�ϱS�6 Y�~���ʀQ��4���@�S�?F(�& ��q,�'��Y�x=n���ߎO��S�uo�F�`�砽/�ɀ:\wN��8�� ����3��S�$}0��e�e�(N�F��D�5:l`�O���bA��+vb��򑻋RIr����3�S6w�E��1)T��(A�TϚ9tJ@�Q�߅�嵓�g�y`��Ё����JX���>�l͊����P$���N`�H�rv�F�b�<c�ϊ%�&.3��T�<��1|b�:�XV���
�d�p�yp�7@@Xɚ��xh�Mv���|��Dt��#>ַ���=�e���-�����ióf��AltŊ��N���N��|��x���&�-@0��$��sh���pO�z�Z�:�Q��ϭ������]�9qA��[Ђ���ۤM�>��wçB�~\�6�ua�ᰰ�]N�Ji��`ԭ[�<CROW��1��]�D�jGt�y�y��qt��bI��t���+��`Gd\V;2*Þ�mn;���ye[�����o���[C��:��Ի����ӿ��
�]��D���ď)_KpJ $aSc��{w˕�OS���f�E�eB�Ō����q��|��y��9�,d2���r�Z�N��Pa�P)Z�?��sbb�
�Fb�8���	ruj]\�GB'��!ș�Be��~��B9�'�^��Օ����>ȹ��.h���ͬt7���-�n^s�sOZ��N����Ƹ>���vr -BtY���v���X�^,/�6lp0�I���� r��~*��!P�V������p�`���G�ߖ�»���>[�r�|�rj�̽H�\�����)|+&�z��Rth�-�H�-+^���><=ʽ�>�ϕvn���a^j����tN�tb� ����0h������N�ѡzI-�:�#ЦP�͹!N�A�sP�s�d�k `/��}l��`ceb��E
{<n߷�[P������|�$�@S�R⎠�E`��(�jwnW��2��֤���I��3��#`�ӳ�Ish�ܙ��>5uh�0�e�	l|
��7�/���:��8�q ���<!��%#�� lq�%�r~!� ��/��и	��\E/�_uR�k�[����%����j��ǦU�����uظ�gj��;�;��VV�,'¶�j��tZw�6g�Z��}�=������]�U�m�W��3�?eߙ�rn����PL��Ч�o[�8Is�R��{��n��=4 Zq���J��p;	5Y��/� �0����%��7��.+�O�rXVf�������&���,���ޭ#\�����N�z�v�L�C�{�-0C�����b�$��H��l�V��`C.�N,�|�{��/9�d>[�ųg����\,�&nW�0�6�͹BUƴ�ʨ�8(��y�B�#�&�yG�q�ЅF���*��,�4�$�UBk=�b�����5��o>��h ��Ƒ��ٹ���'�Y�w��tN���WѤ����p �����r�*x:��n�Ժ�H�9�lB�ۘ�W��� �hO���9T�8ף����O�>ǀ?�:/~�b��7��z�s{���:�)=��A����݅|�9�%m��Tl��*�	���G�E�W�������&�^�%��g�_�!R��pH޴�Tm�vS7e�������׶�����m�H3XmAΩ�{�]�����m��:�'I�~�w�i|k��{=�8Wr�]Q�h֌;yںYG��d�GN�x~ ������5�ߧݷ �7�p��9��g��}O0�)8�?��bB��?��������&	0r��Z�I�Q
B����q�QH)�H�6�����p !�����d�l4�/_����f���Yl��^Q�tÎ��%2�mi�`�_L��o��+i��W���{YP��\+�,�NM[���[ߐ�������Q�'=�Gd��i�S$�ulY������\�J�3��,���]�@d
�ARg�w��ϳ"]�Ϳ��TBlM��ڎ���ϟʊ���x8�,mO֜W;6���d��S;i�b]q�?W�KoߣXAxil;�WD!��=��ʌ�i�Ut���.xr9!ҟ�S�r��jނ�=%&��ԴCF��-�RL/3�tg�'R�4��+����?X�V�`���Z~�H�;Z�t��`L���]�c�R(��-ɩaf4;R���{��Eï��Ggh����W�y���ۤ/S���ImJޜ�kp"~]j;�:cHƘ�f�)�����,��@��Z�r�oЫ)z�H�6���U�X�׹j����QC�]4��H%�̢��'!;xG<؎��C\���}�z���)�pb��m�tӀ�>�[�N���I�Sy��X|_n}|�[�mN��t#�,v"���e�y�x��4v��M���w��6ا�ݾ����ἴ�6?��u�<�r6bc�"����#���e�ښO��j0��V7��Z�Mh
G�*X5��F�n�����=�Q��	l$�3���n�Qw  I3�#�(6���u��k�2,����D!	�� �a��G��1n:(�x�
�X�A�*˲
'7D��|C\\x=k&κ���t��`ݷ~��n���Z9 v�'�;�-��ѷ�g�r5�9�LѾwA�w��7�}7�t�"����io]uO�>uu�ko�U�x
��Cd�#��Dy-:���+�#Y'���߳83�u7]�Y�#Z��������p�Rlc�k��6V�.1�mO�`�*ѵP���r��Q!Ɵۖ�n��m:ؚ�vZ���/�;�k9T�J0�j��ԧ�ˌs�b������G+sR���_-a�^7�n�@Ѡ1d���5��9�CM�Dv#�z�	�En^��TY}��Ӯԑŭʮ�Ҿ�f]�D��E�W�"����fM�X�iS֟�#�c��'��;]<��_��cT&�PG`��J
����؋h�J�08�;�i�6�!��5�~t�
qO���AxW���u�����&��6 ���~�^=b�
q]�N�10%��r�B�S��+��,G����yOۂ�g��q6:'z�t��-?�_V�*�r�C��b9����q[Bi|�?4vc��N�?�T�,������@j$��Q�7Y��؋�p��Ql�C�����F@����w�1��Kʁwh$.0 6KN�	���]��6h�zo����C�n"�%N�Ig�D;�j�-r,PO�mL$Q�耦h��ֵ�k�3�Z�B}����=W&gy���Í�������[��]8�r4z�Y]�݀��_t,d�qGV<�)��<;�bb�'�&�X�D�vQ�H�b�-��z2��4b�T�$X71�Q�t�q�[��DN�|�Y�L�m�,�T[^{��z�B��J�t��j��4|�5�+�s�Y॓.Ps�-i"����oZ8!���՟)������r,wArh���;�v�����L�y�i��� M5�͚JA�(u"�*	l,.0;[�y6P�Ӡ�\*�@��щ��f�ެ)B��3�`*UN�z�=  ���5��)ep��N���v ��RLU���Wuy	��Ƒ�z��.��T��1&�Hhw>cx���1 FU���� ���9c!�LHt2�'��k�����X_������l���ܧ����<��爴`9��ί^�]�C`ֻ��x.p�u[1�:�c�sE�һurHF�]>gf���lls�ה��N}�\��c��ډ���K�`nh��A�(BuA����i�^���=�^�>F��$J��S�ߠ��>ѱ�?6m6�HLt�D�G'*l���zm�(�f�[ǋx��I����N`�H�vu��������c��W��5�-nX���7���ͣ���e��f����НE������Gߗ�U�T��ꁵ��&�%2T�Rؒc�m�KC���ڕ��M�V��Dtb����E�^��l[�<-A8�S�*��^=��t6�֩���!��m�|Cb`@繖e.V*#�����U	lױ�.�m2�GÊ}�0n:�q��62�H��0�F=�Q�D�>S����(��_���A8�I�`�X0@s��N���E�bN�w�Q��y��-�O�YOM�+�r�`&Q5�$�	�cj%v:<��`Fֱ�
J��7qfRa��O�T�~��ގ���e��%����6��=_�Vie�?Q���������pyE+��f����C���R��n7uHFjs
-4�uA8%��nb�h� Y���ն�c<}�9��{�%�P�ݦ�����W���P�Z��8����՘��3uo���M��6��/)����Ӕj�2�N�+6Vzb�`��~���r8�1Ж��Wޕ��`6������ 2��ך�kk�������B.?4N����5�\u��,���k������"�ҏ��Q݌f��Պ�I��q*ҹ���j�:q���Y�f��5��5�r��mܪ7�3gc����ZD"�O��_�P��!4��a:"�-ksCjV��X�>:��#��Ez���e���m3�jx��^��^]���^�J/0r����|N��-o"�r'DcC���d��[H�?A���u��I4ݾd�v�V�{w�<��&�w�/�������5$�~u��Z��.{�}�m߻܅n%��?��jH��0IKyі깾<�1&~<W^;*{rl?ݼB\	��\�kq��m������y)���q�$��M�{���[�MI��m2;�$�n_�b�b��w�L;�,�+#R�Y�G�rΥ�W+�?�^�&vrEj�>]wb���;"�k�ʢ	+�rߥ��:4R0~	�u(�3�6�T���Ы	�1G}���yjF�^=��r� �C	y�h@H	����|�l���S�R>����Ո�q�:@�pS�5�^�����ߗ�\���f?,9������͉��ăf�\���s�H�6��Ѓh��^>�-Q(&��
t�[�N��	݆Gg�O�[+[m��0%��=�2��?��KL��>L7��}�g�z'�H!lCm��6���j9���nC��K����C'i7��u낟�0�z.���L��K�����~k�U7?DZ{%����蔴\m86�h�-o�0��gw�_L�D��L �sCI��ƬQ��j��
T�$͛��{�y�˫kx���7�"S��<���S����_�P�(
�m�~K�hx k�w�lp%-W��0*��=���p8UTl�K��x��#�	l	��l��|��A� �C߿O"����hk@.�񔘶�oh[�F7����D�4$Fݟ)��.}gR��(Ȉ�j��rN�"�a�/7W��'�Ð�C��C�  S�ַk�:��|�^]��c��n$�ǰ 1V��V.����;��$Y�����/��)+���w�.J�4tj���D.Gm�,t��L��A	Z�(eE̬Q`��y�A���5���9t�[��	��#��8J�J�͚/a�Q���p����a��������~� ç��l|�v����cH'e�>z�����zv��9�����<=�5#����c\��e��{�g�ߑ�?��x-F�0�W��!ܠ��	z�D��f�d�g���QT�J4�E�S������(�|��t�є�+cU @����p3H�$L����Fu��v�@�Wk�K�m�-�@q�JW������_�rGN'�q$t_�o��&ݬ��K�$[��rwwCixB���b���N��?���u(��7vJ�Yߚ�}��~���n�~^�ጁ	�s�2VW8t��\�h�٘u`�quv��m��y��h(��.u�����FᥴUiM�[e�G�s$o�Tt���3�o��(R���|�pO�Ǻ"�d]bDAZ���@�7R�
�e1���[_'.�C��Ǆ�];n��!w��k6���@/�����Ɖ&�"�0v����&:����&�q{{K.�i`Ҩ�	��v�S�������؉��H����]J�:B�����sw6�gU����
�3�å�t�2�H�n���]8A���!0���1F�m~l�@"��и
�5?��3�u+��	r�;\��"��̳��Ь�y֊m������u;<�fZ��f��j���ڋ"0��~b��a�(��Ն�E�9H.����p�9��.���%m@���g��l{��@'�q$��j�����U��@Y�g�}_���,C�6*'�vҍ-Se�O�9?�<yZ���lK�0���[+$�����Hf�ӷ쑁MuJ��W��l�n�l�t���Zq�46���%����Av疿�Z�Ƙ�AG�����9�#�N���/��q�ƹVa�F[��ς"-�ab7t�����7��"��\:��z�5Hk�������>�$F)�����e��u&t�1Lf0�D���.Õ0��~�2z5�� =iKU� �m��sx�,SL�ux��e��`��(�񏢒?z�y�n�j��'��WWWp�-�'?�	���ʊ��i�.��Ĵ��ϥ!�ꏁ�p�I|%]` ��i}1x��)�+���w֞��~]�2v#��`ҝ���]6��>���侟P~�����y����Ԇ�& �V$h
�n�I�V7k(�D�7�wT������ OR#�j� ��\�r�w��A�f�E�ĸB' A��5;^��O��2���4)����<����̎����{���K8�>�}���䏁�6?�G?��7��;3~�����5��w�#M�����S�euɞ��c<��!�h|,��n��-�)L��92}>���=6������:U��cA�#���*_Z7��~M��B"��o���d�]S3[��f�Zn�l���<;���j��z�/|�Ih��Ϫ�;��������WU��p�J�mܑ���u0�y���Y?$mtXΊ�U��y(P<Mκ���9��K�u	7��������P��aYl`���j	��uj�q�Q�,��h��D<�V�5�p�ݐ���=K8VJ*�+HIS����f��-�
�k�4�X�7����	l	%��EU���^7�]����Iq}e"���	�^qfh����؆�>��VF���7���cWݺuO����e����Ih��)Uu��Wi~gY�-�����؁��dL�ÿ6T�PY�w[cyw�NN�51>+���j�����s���$%�p6�`�h��;A ��P%��;��]��8z?�`˘ƒX�7�D��8UME�B������JV Fh��B�b�g����)�%�7'�q���6�ΛAE�Y�@�WA�l
��`GV_�*���b�{2��U��1}<
�1�q�$'_���v<�\�M#m�O?#���|�t�u�?r=m�8߅�tz�K2HlK.w��i��H,��.�L@A�]��F�N�s�u״�P��I�r�f�,L$����5�8�pP�?N
���E�b���H�Z����WS��U����2�x�f��Z��q?��s儥�Oܙ`�L[�p��F���Y�A&j��	l	���uQ�3:��a��Q��VF���Yr�N�!S~*�OkS�z]����HSO�GG��l�ޒS���p�`{�0��f�e+�\�mذ���ny�:l׮�~��}v5�2�@dH?��ѿ��O݈4c��/_<�/��ۛ��=mv���pI��)�?����nvG��1#�D�qW8����Q���b�	��j"׹_ʭk�ƅ����'ܤ�^aM_d�x,;�zfS4e4ݤ�d3ض��8��y3[�VdN!�ѽn�����4�ze�����f���aN9�<�!T���!����\��ڸ=���}����b�u$tz�bmܤ��ۡ߷[�n]+ݜ��5��	��D��96�о�)@&V����*5X>Z���љ��mz��~`0GTE�Q��P��9�������[�yXB~v	��T>o�� ePܿ�5��b.sإxm��n��[�icҪ|jSϡ7+������0G����Γ�i���S�]�6��n�w777�j�V'�d��Є��\��@7��
�n|��cя����Ʊ͸���k!��X1�f�=1��<�ߥ��*�デ8��H��9��&V�X��e��=d��w�MAb�����w�)V��R��O��NSrQ^��loo�����'��a�ڲ��7�UH$FJJf�M���eCԿZ;Qr�2��-�E�h�ҡ�=�\�����V����㜯'�q$t5����^^̰D�X��T��8���2��S����W��h�k�q�@n��n�M�ռ���}�V}�`ʶK�nȉ7Ay�-]����]�L!֋觡끲By���n�63����yh�&\�V�OH'%�E�4p��9��)���&��s�u�gz�߂DS�ܔK��I�a��3�l���3x��U��$"�k�ޛ�H�XoPg#%��Z�`R��Lw�=���X�/���ɩ�4A�5�$����b.k����E]�;��J'�q$��R߿z��]��P���%Y���ϳye�Ʊ���̪UZ:&:�*D��l����O�!Y�ᨭO�s�V�^D��Q��M��Th�^w��H½:Q#��e�����M�g��>0�Q�7�`R����He�`e~�]��xY!�V���(p�����CAn�ʴ)!�	�
����J���@�=4O��f`v>����.��0ˮHL�J2�Q�X�zP�WmB�Cbp)S>^/ksϚ�܆��Zi8B:�6`t��ip�'/e5S��>:��#�+��􋟼^�����Y�`l�JAB�\�(k�`���������=ŉZ&��e=n���eE���>����Ѱ����|�s�щݼ���'�Xwc;��5Hm���@'K�Y����e8����7�82��.�A�Y5<&���-_u7ބ����\���Ꮀ.����7dN��2����y�x���>����A��c��}��Q�|MW k����}�*�X7hs�V�5��u�<��\&F��(�����i^T��>�)�������a�R�	�ϵ�a}K�{¡��ge�?������U	���;���U��Κ�JX/�h�ڋ�%Fٮ!-��u�=�+r��u��+#o�[�0B���\�g4]�[�U�*�u��y�|�O����a��w��44�0ϔ�>b鉥�8ڬ��|~~��tO\��9���O_d&�,(+��$��+��4��=cE�ԕA{����:��$��w��-�y�9���������[l�묢�y���OYX���:p����0�]ط)���6b�.����6�u�p�_��ew���R��ͽ6��)�~` Q�2��Sf��V�k��%�܀�o�pt�g��n������J	�e9� (ܤ5r12Z��5�4i���@��31��D(�2��bt7RÉ��l���Nz,�{���?��UQ_;�@�6>��1S�Y�EY\��9M��(E�m69���`��U��iC��� �K�z�Nѭ� �G^�ZV�/�cw�Vޘ�@��x��x~��L'1rc�t�D=����D��}6j�s����{{��~i���Đ1��QH��1(!�V��m�\���3c~gY�`�l��I�Oԇ[�i��+
1���Y�+�GS��9��}��3J�)�P6Yϒ��U@7%�MARRHR�>����w�==7�Dd�l�����pJ���{j�_�BG�dJ�����T��|	Mǹo�`�����_n6�Q�z�����-'*�+�W�-�OH����_�1.ȴ2ӱ�|oSׯk:9��L�����0�e���ϯM1u
���4��}��eE�X=��
M�n���\�K���:�������� �?
X�S�u�a�x������cq~~�l�9�w�RC�h�̚������W7�[H�(���&���8�+�D,O�{�I���Lb��^J:U��T|%!��2̌�Ξ��E] F�Ų5Y�(`k�T,�*6_�G@'1ʑP������Oټ5����&J��t� �͒��hS�����.'���/��SgCs7�6��N�#}�|H4�=yO˿�@w <:����<K!M��M.V��R������Η0x����v�N +��=�����R��iH�k
�9ĺ@� �*eiñ㚊z)�%o@ ���o���.f����Y�֦��͐����?���u9��k�4�,#v��@�X�ԁ)F�M �ƒ�+X6��g����J!��l�ݚ�K�b]�[u��-Y���2b���^�G@'�q$�7���a5G� N<�����%����t�� W��5f��vh�½�Y�c�?��!���8��݄N|��(zZ�Lqw���=��75��fL�NN�%�b�;�h�Kx�2��il�m?^����)\��;چ���'`D��i�����5^����w8S�n�Ql�y�����7������=���=,��{MY�E*@?^=c]���Mި?�ò��9w'yfAI������Tεb2:!����'apB\��)67 ^Cހ#]�?o~'J��9}�6���4/����Xc��ġ��Fd�-���Ԅ�q�T��U�7ޱ�d����^�"�7o���Ώ��{��o#�	�e����>mno��a1������#]j�z8t.�I����!������Ϗ���X�D�SUa�X���F欤XT��5��>�ɇ���s4{�1�E���}́� �T���:�E��ˋ�3Ϯ�ӟ}��_���o��7��|��4�8'j��5C�E��}p$���p��@�^Dfș&eR��?�W��H`A�=�����N�ʬ�	�c�[��C��G��8�g���'�ѨD�$��zx �A���uD��Ŗ�N����1���Cs:b��11�],�6�!��]uSh�t"In�By�~;���C����1�3��-G�8q����sCi��9B4�)�Ӆ��P������:y�r�̿$QѾQF�0�N�d���3D7F�E���yF��6�ճ�����/fP�q����	���0Ғ�I�|�$�)��P[�Ԥ���~�@H"��8��1ފ��"�Fe��m���S�'R��H$�i��5�s��}�N`�Hh]T��b�A$��>���/��Ϳ�?���[�R�����Bx!z
��������8�a���.�;�ᰛ6��MܔT�tb�:m�s�vW�}�.�����7�]ڥ�X�c���vS����7TIWGʏ���C����[{* ۦ��/&�����a�<�!�+yeY�(ʧ-���R}`;n�ݲ|�<�����l���ИqE�~b��$���t�ѕ�W Н���������_-�GY�T?5O��P5�_^���+��8�7߿��g9d����j�|6o@ɚ���;�*��D��t��o�I,r'Tk	��J�^+��#R8`{
2�)���Z����"
A��$C�Ѧ��%d��o��D:��#�T�(fhK}6_��jI����...���9�AŠD���X��k��)}�槛Z�yƨ]�=�-)~��o*�B%}��G�ݔ��m�Nb4|j~\ⲍ�t�~��a#�/֖}�o���� ��3-��! �u��;�I��-�n�g4���eA�)S<�5M`��� ۶2��Ċi�P��8}���j[>r��٠Q���+�[����s�]~g�@n����5I��]�/�je��B�O�UFB��Iǣ$��*�l�/�K�"���|��w��� � B3£y����5��%�o4@"E��b��*���M\��<�Vظk~/�_���Џl�u�(�L��A���������oIc'� ~lD��.z�������/g��B'��Mp��?VF���-y�I�e��h�&G؆�N�����*�h;�,�_L�p��r��y�9HqV?�h`�^�<����:xy��F�##��Fʎ�kGY�p:�����t7����z���OBܷ���Qh= FW��.�K!K9�������{�d-,.��O����ic�
`ۆa��y��q�޼m@�-|��琞_�W��¦�$�������ş@��[�I�P�/��]4��H�N�ܫ�X��J4�N6x�Hi�AN	9���H�9l��(	q'Џ�WCNư�6��pL,�����{��8?h�R�g�=����_~����ڸ�0��ё�f%�i�$*ay���%��ׯ_SB��d�X�"���d�S���c�����>㧕�]N�S��|G��&�6�лr����X�����߆C��I���6��͇���s7��j'n�.Wï��$\ww��B��H�2���ڈ�s�r�6wc�+�~���uR�e�� .��+�͜PB'O�$����o���k'���t�������.�����>���O�3������?�ş���+�����/~_�8�g����w_���O�xؔ����$����yF�jp�Qe���WY>�iZ~�u� ����ڔ�&Q�Ys�Ȳ������YQ��r>��7@#i�l�5�����x��ffY��|�-�
d�����AȆ�oڕ�f�����?���?�W���������)i�of���Z��`CQ|���]�j�Ba?2ͤKRt�0�.�!�qh���D�m6�{�8���|N�W�`�c�6�h��txT���P�)ݖ҅XhG��0�F(����}�G\���o'n���l��q�x��$�������ݶt�!-�Ξ[ϲ��ȥ�����w�K��Յ'Jq��rg� ���b@�q|%��p���Y2c������#J$�} DC>���^|�9���?��������~��'���SXn�f�-�!O�?��뗳g���~����g�gE�p~y��A.�����������;��V�5��V	����g?C��j��a��T����)�*�e�<OϪY�T+�*��<�����mӰ���4y��uӔ�S�M����V:˪3���W�z����ե��)�ͪ��N�${��9M*ԄF�.��4<��
���r�G$G7@�?����E'����k�X�)�c\�}��\��b�@_<5�)	�?u���!�7M�����~�r"�
�v�L��6m\Q��2]�!����������F�"c�Uޔ�\�N�"�b�yൔ�q��~i�I����ep�E\��,7ʢ��∕
��?㟨6bO�l`�.s�-Λ5�%|�ӟ7�gP�
����������ï���'����෿}�j/�%����������C���U����_�J��O�Wp"��8�W�5"q4>���$%!:�%!uT�B�]��D�S�2�w�~&�4� C��7�$�(��u����sy#����o��p�C�G�[��3`��R6��u��B���ݦ�wL�ԍ�2N�<�i}�t�6F�(�J��V6_w�n����m���g\����.�C�u�a\��b..r�M`��.�$�5�+F�uS�R�@�ltߟ�_�S�lP����z�"����Z����|�-�����P9?�����g?��oJ�����'��_��?+���D��8*��f>�kT�uI��p�@�)t�K�rɬR�9H*������OE����/�Av�H�d�r-�/��&RF�����ҝ?�'�.B��&���5����u��{@枴�kC'P�{�=�N�v��q������6�PZ܄�0�V��X�f��Ķ���Z��?t����1��^���a��V�B�@����<��ý������������s\QN����ZԴ\#�IM�i�p�P|�߳$���4(2����I��4�h]»w7p���Ϛ��`~�����,./�Z)��/���
���g���r':(��Ƒ���.Mp�S%�$��� ������j _�h���Q��7���S�_���V<�+�ɻ�L���DI�۫Kba�q�ŗ�7��\Δ���,��j��y+�O�8,R'M�ش�WL���������=m��rjp���t�q?t��mo[�n�>�������X�r����"X��z�[����߉&��gʹ��2�� �g������M�֞2�6�lވ�\[�ޘM����ui9'�/�a�צ=I�{��I�08��G:ڄO�����Tm�9��=E݊G��j%���>S�Z�g�2j�к8o�Fe@x�"F%��U��dMqϯ/�~��V��>{u	�5�]ޮ�Q�o�����_'
 ��;�.tGB�,��ؘ�r���ϚEa	��\�t�4/x�ٌpJx�P�e����E�f���tJ]�S��
�\@C�����e�:��Oq���T�NL�G=ST��ۈp�M��;2N��(x������׿fA�Ӗ�wg��6�V��(�<O������~,�|��	.�A�Y��`�A���8T1R�^�H\,���{�~N>Xsg��C���r�V*�}+�%X���}kR���������_|��ͷ��������ܤ'�qX:��#���]�^�SQ�BV*���+���M�n�8�u�� ���uO�L虮�Tw6���䱨{b�oJ��-!TG�oI�}���x?cb���6�� �C�)[����ϛ���ɛ�1G�=�WUW��nި��
�J�&�-���tj/�h�wT� �"�jND��RA��֩H�0�cE�
�B�[�/hU�5��
���
�9,��&���/�t��D�"�D���8JV���*G��r����[X.��������$P}�@��	LlXe>5�������i|3�ː΅{J�v�p)?,�������<zu��h
�����j(�mˏ��]�˶�k���ǭ��]�M�|����X�����������sl�H����(f���{����m�|�ʫuE����|��[n@��~K������=��Bo��
#_��tGB��ֳ�l��s81���ٖ]y�������gwO3������N�"AؑBal!: �u}���*J���F����#�1��c��A v=t�Xߟ�pB��m�o��>[���=۔��u=�բ�#�r���""5��:�W�@��dћr䍵X�	xS�V�v6����5�-��4��/��9���^\^̒�*�����N`c��j�}簘�
��;_���+NT���?����^h����t�~X������r�������O��<�Z��swW���)cu�D;P,��Y��GO�c:{�b�<��f�{N+'�?���I���i�>�gP�.zFZ�g`��ヅ �(���~6���Hyo��lD�!Ѯ���2t ��l��ԭ(��
��<Ka�Z��7L��p�U�-ׯk�~y���@��
���_V�l^��Ve4�Q��r�Қ�ac]�-:[;3R�h�OqB�?.���!���N�މ+f*9��i��MmJyS��%�� �{0�N�ߞ�g�Ԉmxַ��C�X��z|��De���hMҭs˥��=ʸ3'됑w����hl����GA��[E�Ni�B���wa�I~���Lr�R�no���=+�͚�g�X�����I�.���i( �ÉK�6�h<%�|Q,�慜FįQi
�,�*�D��  ��IDAT�!��6���jb����SP��r ������7/c":ap�d�%#~.t�$q�br�����1�SҦ���}�W�i��֩�<�>��{`������&�Bҏ�J��������:R��C6�-*�5�V�S{�#!w~��w��{e"�튞��
�������)Z��� ��GrF/Qq4#b,���y�s8�A�x�Ə�fˢ,6�B��8q��&�$���|�ꆦ�����60Ks�.���#îS�;y��oY�m�~�݋��˦Cb�w��y���t�-_w����C�b�Z=
��iX�6��g�g���h^#Ch[��?o[��=j_2��$�(� g~��=%5KO��骪��7gVR�1�����|R�D���;���<��3�ڋ�lt2�����z��g�/1w���٨�P*��:>y��G����~>����������������':,��Ƒ�r~�6�I��FՀ	�r�!t�C�ɓ]���cɮ����c2�}h[�qh�ُQ���~9���#�X]O���h�Fd��&���׿нZğ��]}�B�;�X�����f�e�\��=�t'�FF��04�lV���j�$p���	l	U�yVk��?Y�a�]�z�cσ@
��Xà<�ɡ6���Y���w+I|�؎���:5�����oL��x���o�!n��F���ȩ�{��%nȿ�v�NLN��P[�@'O�c�u"�v�e���ֽ?���4�p�'�Sk�*ZC��quy	ϯk��3��֛r-Ѫ�H'�q$�Y�Λ����-����lХ�ƨ��3y�����q�\��)6�hj�uD�)�w�ˉ�E'a�]��q~¢?�Sp_�(����q�����a����-4Ǧ�A]�M虧�l�e>��g�)���6�+�q�(Z��qqq�5���G��q�@�6����&yX-�պ@dE]Y�W�H�K���+�R�v�|�؇��crooQT�rD��&�d�/�:~�G�)��!���r�����:0�/�����~h�G����=FG�}��1N�O��QN�g<R�+�����s�'�w��5����#�����5=+HyJ������������T�y�*]~����6����U�X�YVI�i�n\^_��FBJN��dP�CGAj�đ�Ӿ�/L�1&�~���Z�����u"�s��O'b:MQ�z�CҘN���e|��}tQ�*�:���}~ڻކ��ܔ��=M�����!��*��<P�~���SM�1,��mA�9�`q��K8ѡ�6��&��%��z~���b��3b��d!��Z�E��̒�w�ybq�-���B�$t_�b�^�J����h��6��ƫ�vy	��Y:0�/�!��^}ђ 3���0��1g\�$]�*�P��٘R��`c(5�C{"?M(���\�W�pH�_�꿰EKBb�Y��� X�Kz�Jh�v>_��L{~q^���N��8*ʪ��y���Xo������7ߐ;����Aҧ�j�T����*����!�������E(��D� �h�' �[�},�U'�=Y~H��1�PZw�>D�b���]��'����)㛧�D��Z��g{u���-������>����X��d3&ǒ�b���O��M�lN殘�/���Vkt�U���N`��tGBU�wY�(��	ܽ}O&[��s� h��5�Z�rG3a!k�l=<c�m���
_�ܖ'�4�'�];%��qH�-�p���Kt�;�ÛE�.hh��'�n�{<����I6�:�)n�/S6��`��P%3�wﴯ��_��������_��s���������&�x���§*�ގ���UB��p$��8�$�G���RO�#��ς1�~-����|�AGl�SJ3����T��kL�%��es����c��&e
��UB����zQ5i�z�ޜ�Ɓ�6����M�)Wy�L
�:YF����W ��Eye6a󙥤�Q7�c�����p���*c:	�f�����"[3� �_8��A��!u:b���z�'�����g��{�4�=��S�n��������"A	��lzv`~oۧ1]���Sc4X�����w=�#p9�Y�B��2^��۷����a��P 8�&�}�~|2�#��8Z5�Ue���;�Ϟ=�(�����u�:r�.x@��`��]>��-����z�@�>�i�v�s9V�H�س�Mce�[�C=��=�r憸D!ݦ>y�>����:n.�l�xW��>�gR��0�t"��]��.��4���J^EU�4��xC�;*���;x���?|��7�Nz$TW���*v֥,�J����$) ��#E"F�-LC��X%��֫c_D���Q��	m��?���:	S�D�7�`��c��J���6��������+f�xYĘH�Ā�<D)��c��WC�k��DL��v���X�S�q�q�Dq4�P�J��-�쪹~A��b4���"��N`�H�"����y����{(:��U�\�6��Ւ�;�L��d�����Z�)��8�*R��S��9�n�}��^s܌�G���b������>_�S6�J{�c�$^�c���@w���A�X��j.O��w���b��R�^$�� y	l�N���YFA�(��
�n!�xq���O�_��)�I_#D��Q:��#��/���/���6�n��@�Jj��g��)�f� c#U1�ǥ����{L�ߦ��G��P�c��u������J����mܦ���߱��b
�N�(��trZ�[s��-�uǿ���o�1��)����##�s�� ���?��N�Ptl��5����װ*V0�WP59\s�o���՛9О��6����<M�fY��|�Һ.��l�o4��y^����b3�����b�ݦ�F��B�{�=�N�v4�����X�C��b���A�f��O���ƸH&ȟp������O��9��O�D�3S��E��n$!`;�tʱ�'�)�a튝�`ȓ$U$�&ͽO>��,c���W��w��˫+��,Y�'1ʁ�6������˪��裿�y" ��B�ˁ�	9�D��ï�)e�C��>.�'��N�t���b�쪳0U��o�o+���{������ga���G�ѹ��-��.�='iw�?�^Ԯ8e��7؏�o�h�}.gc,��\FY3��u	I��(�<��
x�<�����My@gs� �*���X��J'�q$�l��ʲ����(4{}�7oސ����9$ ��R���0��'�L�c
h����z��-�|����|;���0v�����;a����p��S[H�-ؾ���G����ꁓ�!�H���uqv��B���Ƣ�m�Ce��Dm�CvL�-�Ncy�,v}n�sz��0��M(M���w�B\����D�<wu���^�b1q��(�n���zӀM�j�f��O��O?����[H�r�Bu&{�}�� �.�j��I0XF"�����4�Y��08iPQ�0;p�Te�m��<�vlQ��oK��P6��Y���}ܺ��},�B[���5t�T�@Z���g�p��h,�Jc�?mlΌ�!|�8hi���m�`'j���\o�rxi�U�jҤ�C�W�mY�5�c�|���c��l�.��I�r`"�q������o�Kp"�x�Aٟ���L��D�A4Is
�	�$�4� ���]�]�v����e������i����Ci���R�;=�ʮ�������xf��o~FLa��������]��u��m��B#��l�w��@04em��t���YGQ4�\ ����P%�����aI�]y���I�[�v���HHm�
�l�f3��I�|��C%+tP\�]��V�Z�o��a�FA���p\L��!��P:�.�`"@�l�Ѵ!C g�}���*�E�aJ�m�0!�. oh�������X�\��_��D���{Q��bݓ8��:�9����JҬ�Q[G	��-Or�����X���u}}����G@'�q$��_�{���E&�]�3
71�ICʢ6'�S2�>�I�[N˲>�0��qbeӢ�cmx�Vj��7�f�a����D���x�ޕ�' �>Y��aږ�f���W��p��($�mu !~�ޱ����4Fv%@�H,=�gd��5��kU��IfiFU�k��R���	l5hz��98iH|����Qf|�	ׇ��Mĕ��Н�Ҹ�����El4E�rH�?�,�6�~����Iu��n虩�MI;��8c�'��Q�����qDB4�K2�{2��/���#�j�HM�ŔJ)�|��`�,���-�(*������Wp��{T"M�=�?9�:0��Ƒ��b~yqq������	�
���a��2@����r[�cQL����B8�@i~�ï����a�o�@:u��^�pMQ�=$����o�&��W_W�3�A�vܤi�6�P�ڏB��u����b�`jG���4�k��Y�`t6 dQ��i�aH�
]�pR=0��Ƒ�z��Flg�jI��'����}��f��G
�F���&Mj�&�� .�bl�Щi�d<T����8���5��:S7�!ݐǤP��N��o�ƀ�6:�|����3ce�#�ݐ�11ZL�oM���⿷?�S�����vvVqX4�ELQUPR=�g@����{����eUm����<Y �A�	l	U�M�w���O��.u	�w7�Q�Y���P�]9��d֨F_��M��F��蛋�LܲQ��+�~�R�� ��f���L�B�=����MA0v*�%q�[�I�_����]���k�>
n&������b|��������f�T��<���>��6��N���vd��֤�&�-G0\'�w��e���`�f�kI���F�זk�k�P}���{�̫￷m �(P�q�Qީ��Q���;$�2lq'λ��;�4+�K=p�+�����r(�,f3�RM���/.�7�7�[xv~�<u^��.aG:�0��ƑЬ���ź�	C����f��'���6`��`���	9�8
hO������,tO�]���\ڕ2U��oV��:�A�<bu�=���F|q�p���8��<��ُ��/L�E}��d�6�Xږ���!tV�����wܶ��tT�Y��fyF�v�Y6��b� d_�����������J�d����;����6����b�\fh��V(h����;r��x"i����h� }]�),�1:&�{���:�v��������DC�3%G�~��~��Ӯb�]������_�1Q���!qM�y��Ց�/�Em�P��Ձ� �4؅^����i�����y����"U
u�NtX:��#��o��u�g8yУ��G�i-@�L+�($�
��d��IS�_̇��o��7�X��L��җ���N��{�ߖ�?�e=V���{�}�:�w������߆��<�鏶'��8@�6_��,e1Z�ՊA�1�JEqe�����A�S��r8�A�6���4��,K8�Z
����ETȟ��� ��=5�s�Պ$�\��&W<�U}�a�l�C,� ��,�� ���0"F�w�߅3��s[���Z�K�K�s��$+ .�D�1t���s(�[�9����_Rp�o߼�r4��ֺ~Z��?:��#���g�fBT�MI� ��(����ߠF&���2}��p��c��A9�v����{�EM��Ҍ��%�=R�(=���01t��U�c����	���=!.�V�{d�;T�d����9�)����(([�Ƣˢ4���V%���Hr�D':(��7�����hP���k�L@v�����0Բ\��{ڇU�H�#UwِV�`sՔD��،�w��s��?F���K��7�%s������{2���/��_���1޸�9C�C�v}��1Y8��đ^���Is�����fMYX���E��|�9<� �~�t�/�Nb��Q��+�@�k؜�-4N �l �@�^����[��!��X���d[Q��z��	�1e��F&=�Y�7��x���8��O��ʁc�f�
�����C�*Ly�S�q+�� ���ehM�㇉ǡ��1tf��#�a�\�N��n���<����B٢X�C����[���3����o�U'�cM�-��1�*Y�fb�d��.ɧ����\\\�ruG����*%I�.��ߗ�*4es{njݴu�^Oi����2�ӉbJ.���W�M�[�6�)���7?�h��U0i3�����"��נ�/�^��e��|0�O���tv�'��"4(�RN/����_��gc`����Ms�wc��ڣ<�c��]9��9wLE��y�H.$�P�Z����ʊ�B�1���*
 �!����7��5[�5}�3�,=���6������^����X�)jM��'i 
�Vc��oMa�+�'��>�p��(��<n��S��O������y���q��J3�}A�	44���g
M�u=�qi���x�����ъͺr3��]ѡ��*���e���QbR��d6���~�%�?��7�~X��|���l���Ɓ�6��n��f3�Qz~F�BB�#�@�~�&����l�Ǝ-�S�c=H���,�UL��>!�i16!��EgW+��h[��]��>d�n��\��gv�Q����ڻ�s�k/�t�C�#��pR�}���rT/gt|�^4���p��'�I��̭��(�k�BUW�f�- Y�#��Ev�Z��ƁiO��eOHjp3^�qTf�/�:I2��7�k�}��&�B�&%�ɳ�t_����C�{��?���N-�ϳ����?D�C"�ts�I�m*C����}~����%�~:?�����ߖ�83�ѷ�������H�(��T��e��犔D/��м����V�v��iO�q<{��4��k�L�������jӠ�� U�{u7
�N�c��'����V��D;&UCP�X��Q?B��yt�"k?f���;G7㏣�4�}:4��ov�PEQ�͡
Ǉ��qRp�j=_���s8;CN�R7�r��������]���$F9Z$gu���(.����?�����I��R���k��R�>�9�������e{E�}hLWa�Lх8T�1ѡ�n��>V����Hcb�Ǧ���C�R�=�Э�˞;P!�B����ǝ�Fl*� 6nnn�^={�|{�,��?8?2:��#��Z͛ɑ��aڱ��e��@B�lٟ��L\7�������{_ڇ�cǺ��Ã�.�R�W)V�S���8I�:	O"&Nߎ�� RfJ��Pln����y��w���WnF괟E�f]���=\�J�+������r����Y�zy��84Mǣ��C%��M*j0JL��޽���d��Yj����Ҙ��n@�]hp�:z�S�L۲����p�,���F�P읿��m�����	pݥ}��*Rg�����C��àS =M�m��V���v\w=l��u��c��6���G�e�q7Pἦ1��<�r�f�m�U*Pɾ��9�����o�{�|v/Ws�<�hN����>��&���xl�
��Y^�%�P�8?�lfcJ��[n�iB(=�3�8��v��߇�ŷ9}�����~������翮�a�tg1�E��?M����C谣�n]���l����QR���l��ء�]څ�3��ۇ]���Y7��<�C��!6{��	9�v��Yս��ֽ����g��J����WP.��##��r�6�#]�6/�g#B�E*&�`m��KK��~�c�̯1�Qg.t��8��܁�x�@j"BI4�������r�����f	y:��,�J�����a���b���YV�뇓�Ɓ�$F9�i�����j�����q�D�4��d9-"2%Q|�nw3��'<ʹé�X�� ������[��j�	r$M���?���A�����S��]p�K?���6,�N��ׯ�P�!:�(g�$�1}0g�a'Vu�ܓ�֑vnxC�JO�{��cpf�9b�͂��/��f}MrD�S5��+�/�a��6%b�*����NtP������~L��\U�N�ʫ��b�6��f<Q�I$��'�6�����Т�*{My>t2�x���}=|��c�v�����A͠�kBB���rc�L���=�S �ӹ�q��8�����>����q�hv�1��w�o#�)4��yL(���Ey�˲�*��R��t�W�pu}����\$��Hյ��D�(�8���ϟ%�D�h.hp𣜑'AB"��*�4Wk7�h�:�#D�"Z`�N>�	m8�)Ş��rɭKLn-�����ym˹8T�{��I���ce���a�O�?T�%(:�C����d��8�o3���8��2��d�p�F�c`i�f_E�*ۓ�D���q6o��Ni�=�a�$F9�Y1�eN���ik��P�X6 #I�U]���`�����c�4e!��i
�g(�!�z�,�\��㘮ʾ��gI�u��'z�:����?�^G����S��7������Sc:QS��_���4M\i!��۫��}@���,���= 7�Y{����-Vf���:Y��>J��C�\䙞����B���2�΍����'l<��)N�~�Q^�U�2t�г��\��c:���Ƴ/�H�U"ܤý�����|W���R�Y�nMO��co��)��^���`۟10��7��^�#���]�VkfҌF&�Eff-��]!�[U�0I&��C��?��Ҧ��z7����{]����/���������6��T��{>*j�Y��b]6�FW���<y��WoV�cY/�#8�Q�g	6�_������E��h�(�d��ꫯ`:��.����f����îF��x�Bߍ�?ۡC4�>�N�z�t�N͆*�f�}̷��ň� �>Y2�ىw�+ �b������>Zvl���t�j)t\����gU�v�h��4�}����W��z,$uٚ�w�ս�[�|�]���������h���ժ��X<P&�$��e�^\����L�wd�»׋%��jg:*�,�Ʃ�>�����l�Z��'��g���O>!�� �z� J�6�<MK���Ʊ��Z�2�^�k��5fՈ�Ol1��4[.P��KC}@�K3�9�>T��Z\���.�y���9��d	��o�?'�a�����"��s�����_�r{wC�z�[n�e�P�6Bc�ꍠK3�^�F ��j�k��w��x�<���gڢ3�x�����p��2c7a����n�����zu�z̀#O�6���N�1(&�Cԧ7����Z��v�_P�6yO�y!F�gɈ��#Mvw�ZW@�c������;���*�s+�FC��5�l���냭{�`:vwg�Ү���I.�p�q)7���Ƴ?��eI�I�ԃ���9��.�l�%��c1`P��{��*�����[�a� ֿ.d��㵶a�<[�a�FI1o�*Y��*���[ڌ��hK�4������t'Bo���,������w����~K[ʻP��6̫ͨ�4bL��9��Wv)�O0�
.��+o�K�e�}P_���|f�^�V���H�����>���BS{� �ݺ��<�m�=�O�)����j����0�3b�c� K���ں�k'2ͫ��
�<�������~ ��l6����tgC<��tH������o���MY�D��:���0V��
z��t�ҏL>S;�.Է�U=r���t(3Oz�G���X�z�efh�B[�"n�����@Y��gcynx�&�\+��v��>R�X:|��iHp�-����<���I��������O02�����q
��>7��b:�q��Qʼ5'��>��#�l ��@��ӧ����ߔ���J�gϟ�_8��D��/eNG�cǲ�h�kBh#9LHř�p!xH�c����Af{��;2s�tN��q�K#�r����_�█���9|�*}�����q(8���Z���صnc.�.ptchn��"B�#��Oh�Y�ib ����U�ۨ�`2×_~�n�o� M���Mu��q&Kg�q"��������8ip_L`��R K 3`�8
�D�ƏK`K}�M���>�.q��?�b���X����g�w�|Hu_�}r��ń�c��jjP��W�h��/.��J����
�nz��h���ۍQ��˯�Kq�n��\,�`#�����S?�����$���a�R0�'UQ�{�M/�rd�yz��ud:�����jI'��7o��n�[1b�HF�G�m���V��;&�)Ůyl�q�߿��}ԥ��1Rpe�!m�4���2�B�t�E�l�4�>+^��U"�j+����0��|����'n!p۰���/�˚�E��a����]K��<���E���졵�����[:yy	��Ǯ�"�����`�D�2�Xe�\_=��l����-��s0PO!tN���V�Iv2�w�"�weF]�vua��0����_8ڷ�]����h���嚖+K�7�׷�|�A����O{�кs���nb#�]I�G����y`���� �Ɲ`-:��o[8zˊX7��I�.5c�1�������)BV�`$)�E1r�8~�kJ���(Ǧ3�8�_.���<Y,V��e���ŋf6|�ZP���/+���u�e)&�Ǜ1&�<��l�U�2¨�<��x�
i���`j��g��,3I ��>k������_2в��Khsc5��}`�o.��C\%
�ࢮ���G`�!�<��w�u���"�|�,8��M蛿C-+u=���1�Q̒�x($����G�"�F�����;�xn�\]�Jg�q"������7��:�&py���W ���R�%��P�V��qz�V�u����h[�Xl���? ��&�{O̜�/�ښ���U�L���&M0��Qe�fe��K���v�?��?Dx������w�.°���^ץ}qM��ۤ%����z���q��
:��/������X�:��vg��#}�8{�(h�j��n��������R_#�HTpL��gc6�����N��*Fe�O�`�keeK�ؖrp��)�H���W�]�sj�|s>�ǆ�����7%�����0�^��EO�<���{H���c��-���^���Jg�q"����@�i�+V$:_, V+�L&�W�ͱ��l�9�N�L�ZGL�Z���ct����RdJg�.�i1���p�R����i��u�.�$���l�K�w�s[�~+��q���U��!V��AKxE�,]�� ý��.A���"�}����:�C����5�i$��A��Jf^&E����� ))6.O5TŒ3������؎Lg�q*�#s*V+3��������=i]h�۬�b7&��H�uѺA��Iƨ�ѧE�Cq�'�A���vWG0���(�]����*_w�6��H �����j��q��+W,W��p�����u*���]�'����Z�9���������﷫��C(�C�q}�p�FyC^�S�Q�.���,asW��ׯ�����@�n=��x<U�\S�_�^\?��Ɖ��l�a6�T���|�ј>�k��7��Nq�]��~s�Ґe}��x��ŭ�����)��Řo�)j98�+�}?���>p:��w��;��{���.�����o�=w�.�����f�m��:�c2v���E��}��}����P{�׵��A���v]K��Qb:�r�� �C��l��=�Dnc:��=L�3�@�Ht'Bף�;��lWח������<�N]�)��(�`n@�k��ny8b�PM��y�,����ξ�
����C}#uh�ӯw_�@�^�o`���j����ch������:Dl���%��3
ܶ��c.�`���r�t����־֧.��$n&?X��)!^p���5Ǉ�Y�w�J��>A�F�|�bsJHm�bS ��ϟÿ����{xx �Z�D�Mg�q*4)��*�r��|�����捁 G���5��t
j4����c<�p
:����0ch�q�=���2��tT�t�@��1sm	mf�)�c�$�ݿ't��Z�u�>�K��6ny�]���>u�y�sB�z-^��>�{F��� �Y-vC�x����U9��60i[��8�q��p�kH䚞LȪ!�_\\�J���t'B��<�������?ܛS�d��^�dI+��(�%�����m3��d�2���ԗ���W��DM�G�c��/ǇP�n��
��w����zJn��#�]��\Ȍ��V�􀄾���<���کGh�T~}� �ky�[�ܱ���Eh\&MYm@�J�ܜCkq��v'��	��z\�WP��Oᯖ&�#�l�-�EZ��0��wH��P�qL��wsX�V�)�i;
�1�>C�i�!��W��t��,�@�L���g�Z�|1l��.���cRh<t�o��q_���O=[Z��^�&x��ɹg�?�v��oߥ�xF�@��,T�X�쑭k���C.��κ�XRv�,������?�gv�l������w��F㜬d�0h��DpP�D�wwwF2~���Zz�t'BWO���l��>}
����(�-y-
NQnw��-#[��-h&���H��:E�B0`c�]`�����<�U����ep��mT�u��C�����������w���>��UG����Z}��_���k��t��yX�=�.����u�)�4T^ֺ�/��Ʒ2b�q��P�Bu�)������.e0 �s�t->I���DW��h(��*�)�^eP���u<���hݨTAVe�36?�&��]]^��Jg�q"���h2%����f�td�˵
�HHqB�$��U���[��cϝ��Z;��m1��f(;��`��C�:���%���P�}��l?���ChX��Ҹ}��rye�ڧ�%��*�O_�n���wϹ�HZ�,��2c����u_?����}���kHi :��4

�!L���ٔ����W�M�SNUn�G+GY��FlG�3�8*����"�	�����"�$�ǔ�<Ix�a�&���QL�U�Q�n�:NG�Ŵ���j�p�16.x}�¬��`�:��.f⮲C��=�1F�
����]�|��tî�պ��n��W����&�cB���>�޽2��VE�ב�u��oː6�h��Z^��󟳨�ol�@��&8�E��������܋���tT:����zcfD���y��j�ALY��501�aL�J�Y�h�8�~,��׼�O�c��L���i��:���z��>���jQ���c��!.���w�C���-��CO�C� ��z_]V��s]wLSgL�����=��t�c[��v}��������u���R�JM{J��WQ�����-��q���)G��g:���t:���2Ap���_�d2��rC�>��;��@Ѹn�*����#Y4b�z�e��M�ͧ�﾿�̈���������x�}a���	�;��ϲ����4Ҿ
XÅ��SHh��^c���/��_d�w�=&�@��XDB��.�E�[(t�X�2�~�M\���6#�,:Π�ۃqx])�q�a7��gp���l�M�\?<,T6�W_}Ϟ=c�IY����|m�����c	��eA΅���-{H=b�랾�(�R���Ϻs	��:�&d8�j7�1�i��[��'�}��>����(�(d��j��A�Rfq�Ѻ/�V��o9�=+$�ݶ�ǻ �
���V^
67 Y7�4G4��85�QC�0�?�
�rT��p��tT:���������VQ��3ic '-���UJD�2-]E�cQ�v�e���%f��蝘[�dm�Wz����*��5X8�iǀ�1����o����C�8�{C�<4�rB`9��q߲�8�qW�>KK���F���ȿ6t�1�{��4s��X��"k��]����/��36t���iv=2��Ɖ���^_���%����
~�)�&c*�	�h�`�(M���E����jң���)���HsYp�l�~m�M��=^�cP@�b�]�q�w�y�	��P��sh��[~cىk�xM���4�t��ڷ���g�wӈ��o�賌��e�լ�������@M������oS��ce��.�j�e�)�)�J�j7M ����n)[3f�]?�wo��\F��LG�3�8�Y�%y��hx{sK]��� �9L�cZ޺X��K*Oa�����uםlV`�*4: F�?�kN�ך*+�C��������)���K�㕗CC��њ���rW�����Ä)�{b�݀���[C�	�X�]�c��٭�*���o��v�<6�_h}oL�C�����r������i�����"�U���(��:�v]}�g�QIF3�֨�OS��u+OI�ƶ8 �>� 	���{�ơ}>`�gy;O��ހ�v;�@�b &4nR���I�`8�^ޚ�}�n�"7
\���(�����n`1_Y��
x5���ؙ�t'B��ߌ��e�C/.�a2��CQ�f�|f����fFm`i&ir%�z޵𘮔��ҥ��EJbN���E�u����n�>]&��=}����U�w������)�$�����N�����^�l�L7x7T�k�Շ,#�}M�b�kA��}C��o͑�b��>WJ�Y��w�8>�.7i���,7�eeUBn�����UY�9K���5��t'B�$���i�֊�x\ow���d)����l
Z�����8���2��E�a�x�U1]�0d��)hƭm�`�g�C�N_����]sH��}} ��_��!��^�'�F�3�Z__���{b���0D���X�B$�%ޘr���bc0,bu������C�thNق�_��߃��8FÀ��a
s-��3 Q�9f��t'B��|q{}yUTE��%'����O>���X�߁.8!�RJ�]��u�_���xL�P�m�y�S�U���e9����]?; �vqQt]c��_׻��z�+H�z9�Pu�͘����B�{@xwY\p㟓��������wh�7t��=Rho�И�均�Lv��(hlʣU{)��$�W����<��Y|R��l����#�l��6eah��_�XoȪ����˗ �������2�( ��T
�B�t��∙K}&�e^ݳ�5� X]�yھc��3��y}����b���2d㬾��2�X^Bm����.������P9հ1��w]7�R����t\7���w�}@z�\4��l`���f���y6���\�u�"�|g:*��ƩPQ�f�T���0�ݫW�`�\�^)�߿�I1�d�d7�5�yګ��:�ik}��C4o9{�7�!4���FU}�p�٧��r�@�z~�{�/{K���\�P�[���4o�Oe��?Vf��r�"V��\�+k0{��o}"|)h�}�l �r������E6��,��(?�Q�Lg�q"�t96?�M��<yB�q��f���t��&-�J�Mcn@G��yx�	��ɵu�U�Tԍ^��κ��~�ˮ凟�N�ԡK �j���C�/$�@J@��ߪ��6ѻ�[s�*�q�P} ��b��h`�)�+�]�׍~+�2��]��+/T�. ��<���~�MN�%���z!�c�8��'�Sk7KU=�3����2�3s<�������Vh�@t}uu_|�9��h�  Y/��� �8�c;w��c[K�Lڽ�Z�ஹyW��U�P�in�p��!�҇��?D������?�~	]�H���탍P�|�v�w�!��~{�������t�o���>��*f=	��ꢷ=)4oB�W�l[}t]?��qn�
D����W�L`v��,�ܭo1��<�3i��t'BE�I'өF����kx��SF٫���T������h�GX�����`�^���Xŉ@��u�q;D(���P]���.n�}�!-����[�}~={�|�˻��w9h�Œb����=������-�r�ӫ^��VY[m����~t����GK2�nũ���ۯ}�ӽ�}�[֟�8��ߢ���*>>p�M{���q�D�-����OW��7b[,����6WWx��n*�WB��6N�f�˪,�ۛ�5�z�z,�WT3J��/�L}���g\a`�S}�F~l7E_�}Zސ2���wMHhŞٺ��𝟯�o�ϱ�b�����Xb��69�'o���tYTb��^F�P��66�Y�v}7B�����y�P��KHt��I6J��L�k9�����de��d/^����%���8C�L�ɀ�A�P䅄������iK~�~gš&���G���n��_~nԧq������{��ٲ�`�����o���x�@` 
��(���Gu;QZ�=RG���\c�1����<3%fC��I�^�t���t:}g:*��Ɖ�� .��^�ȿ�������>e��MJ�9�3��S��4P�_Mq���>-�g�]n����hv]���C��}�*����s�XMv���	�̆�'�6	��b��(ny�����.��C�A��>P��\L��(i����Ō��F��m毮��`��t'B����z}����͊v%č�X��%��>j�ɧ�@b�m�[.*�8~���b��/��/�b����2Ѣ�P���;�_L�F�*��.Qk۪��W߾:yr�m���]uu��ҥ��9��+}A������b���
����t'C�j�^�h���0����Ph��7S�������ԧIm3�n�w���Z��¤��r��k�~i��:t��w}�.�|��sn^k�Hg� ,]½.;�1��tu���J]ׇ��u}��=�H�.�(dVI�=��h6��ﷷ �ٲa�ኔ�r�8�Q�6N�����fSt�Mg3�!-����o�Q=�U�gP��@���*x>|b�v���	�=6����ij_�m��w]�c�^���P�����G�#� �.�Q�z�:�VE@S�m�;t,�j���ֳ����Ɩ��q��Y\�"e )�y6�Mg�q"��Y1�d��'O��Ϟ�(�����I���Y��L�M��
'�<>^�h�w����4��.1	>3��U���>>�P���޵��ݺ���	����.T��aeq��kܾ��5X�,+�>�$�/c��}�1�K�;l|ǟ!<Qo�<]�!��o-��>�8���t������Jg�q"�L�\���qAa������ �ܼ�
R��ZS܆2�sX�>�GVV�&�ڳ&��e����bv.�z��9�ǭ�u�����
k�t� 3R[� ��itT���q��5�]5�]��	�]Mخ��/�˿�?��L[��CP���� �D������32N��������jY&�l��.���Z��ux�5�|S���c1��"��иq�!�=�?w~���t�T�s�=��w黗B�Q*�%���C�$ ]�gc��J4��$��)��(}yi��f�p}}�y��3R�Z���Jg�q"d����jVF0cR�K4��X�'vbkb|2��$ȅ���E.3s�F���{O��.�bN�s��w�1�ġ:�	�{��+s�f�C߅���B����c���}!0�*/p����sG�C��Ϫ�F$A�S��+�oL�g������N7V^���{�Ud���Uf����bÁ�h�@�ޔ����_/��Ɖ��r�!��7`������l��(isTZ��A�dJ���o:}\ ��E!�̪�>1�T�Y�쿋��Ώ���Ŭ�����?!�J�V.��U��'�q�u���.@z���&P�}v���b���MG�d��W���&5��_�E����Ϲ���np(�-q�m�f X����.W�+8�Q�6N�r�]�������/�X� �X��3)6��Ԗ���%T3�\m\/�v�L�]f��}��p~Ǵ�c�m��^3� f�v��;f����������>���]�!������F�@�v����K�Z�*4Һ�W��(V>�0�Bu�}?�UY��]�վ���9\��z���Cπ�'p���l�eU&I�0{��_����,��A��z*]�������I��ߛ���g�x+?|Sq�Y��c{;�q��S�1#�M2��]��?v��R�?u��)&#W�Ӿ�e���> ������.��*����2Q���|�c�qI@�\'v�OPT/�Q[#�0�`B/�CŎ��]!W��ۑ�6N�t���F=��Û7o��_N9c���XF��M��&�����M��uʽ�E�.��،.����c_����r��x�vW��Ӎ����	�^�S��`�ŭ�]G�)ڸ<?6��ې���廫T��7i
ާa�q�K���9�F�=��R�����F�qi3�*��E	���t\:����b�޽�W�^�����>AJ���eFu�o�c�IE��BB�#Y8�.�C�e��&Q�x|�_T#11�P�1�c	��.���f����٧`!9��}��!���V�e�rPi�@�Y�I�=6	�˯�.��� 9o��8���GC����>b+F�7��l�h�0}N+O��f��2�ө�kM���+������J[`#l�:�c�� K3�Ǹ����N4���iK���7O�fC!1���s_�s]���5�����a��|�����p��ul
i���D����_����y�:BC���J�վ.��U����׾����O~�c��@�r��l���w|k�O�1d}���t�8�@���A�F�i���Bf�\�����(Ǧ-�q?%y�����L&�/_�l���M�n e��jk�l1_nMh�,Z�'�>~�6�l�����ʹ�Q���j_p������3-?"�����o4�]f�o���:�}19��K��T���xq��W_0q5��.7EH��)_���k���=&B�����e9�����Q�ݱ��m����>7O�E��S��:6C�7��-rG}�o��(Cߏ�.	�R�T3��\��6J\N�[�`c2�(�#8��t��('Bϯ��/~��ͫ`c�5FD�4��]%����"%��4�es#���"��w�Đ��u����ر=�-o��w)���]@�>u��|����]����PLغ����ʍQW]��{~��,5���>:�e��:Q���%Z��/IrH7%�L$Uy��ze���<Ǧ^��9������4Ϯ�>�.W+����g�ؘ�a�F�2�(0S�u�$iBQ�H�f��Z8�F�M�sp��G��/�˞|m�e��c�Z��M>6����>m�����U�۷�]�X�)bm�py~�����f_`,둼�T7֝ �N�a<F���7���^,�]�<�"~����LG�^�q��*�2������^<)h�AY'N������ǈ�%���E
��{5p�5Ҝ׏"�>�0����p�S��n��������B��êk����]� �c����O@��)�w��n����Ab���=�ׅV���{�9.qpZ�)Cs>�a:Ë����
�
6�{#8�Q��F9Z����.K�&�)e�{��=nж�w����E	c4��1�d�K�gj���S()T,�⧠>3�7��s�"�\7Uȅ�U�!.��up��t����`:�f
	��u���+;�B\��-~����Ž�O�>`�[U�~4�A����儼~"����Wʑ��`�Dh�X�p�+n�����x�����E���?S2r��j������S&�e�:�:��!��:$&a�V��=���va�����.e���Y2H���1$�E ����=vL��R��c߸�!`�o��Uh.����������W�``�-�CSǍ��|����h��c���tC�����9�ב�6>2�H�������&�l6��gh�{�����u��}��|�w��]O-���zL��er��Tn�����2D0l1`�8�S[4����Rh�x��Ӑ	���ҽ����8TX�YIvuW��q���)C�R����}[�2�	f4)w�~��|���r��}	뇹���l��`�#S,��64�W�x��5\�.(��z��b��+hf�U�0�lz��f�{,�!�@ͮ�����,+M۶���IC73�X�r��Y��CZ]H��|�����׹��Х�m+�
Ze������7]���/�w�cƶ��/_p�.Ȯ�v�)voߘq�Ũ��cc�=�Ɗ�Y%ܶľ��gh����_�`R��Lo����� �5��V�K��S������͇w�xx��Ԁ����jǊ�8O/ܛ�`�D(OG0�.6p��-<<� S�c��gO��|�A��âx�J�J�4A�	���j�G{b5�f��Z�M�ͳ�"�qbf.r������Ή�o17��U2�&U�+��(3Ox�q�p�N��a�]��X�^�p���^a�4b@ ��	��{O}����%|��p�y7�S|�6��q ����mA_M²<`ͩ��n
Px�ޱ_o	@��;Z������Υ��]�7@��+h�7�� �RpC�A��8���rv5���޼y��;��	�y��
��������l�=�����hT^L��o��^�`+^U�Z-͋*k�r��M:���)����X.{�<�!�g�Ց�%�h�u-���$�e��V����]�������w�Ğ!���x��!��u���]ʋͯ!֨]���<�k����Chՠw��e��� �D��s��9�$_���4�s�98�T	n7?����Jg�q� �|������ً�0���*1�e��Xa�`]3yt%̠]���'��&xl1��}�W�1f�������3_�[~���f�!C�h�u�c��@H����7��}�]�[[��H Q��
w鿟����Ѷ� �p�
NS�1�5���r=^3�L
8�Q�6N�4,W����uAI��p�Lw.(������O��֋1��B�e:���\��|��iO�BZ`��<vm�� ��.�i�!�K�nv��n�>�C�j���A�h�e�X���8B��cXG�����u�_[WK�h�ݦ�ݨ��\��7���T�����%\?���0��E�)�O��_@r͓�пf�ϗS3���|��7i�xD>i��8MyUq�hZ%��wvL2�
�t�Ƙc�#�N�k�d�����9ף\a�[�z[p��{�����e�p��f�&C�=�j�zw�l��"}���e�{�x��5h�w7��1,o�M�c��eYA�q�g��z1'p�YC��o�uc�^��H�$�<������k�����e������O��(��{�ʜ��8�v��lC�"�^� �(���{v� �*oP9*���Ҿc�s�b��'f�?��C��C�z(����{���^�U�C��|jWi�^)ײ���H�r�RҦ����+x��)uO�<�M1a�Z���?������_�ϖA:��`�D��
�*6�;���7�1|�Mi�MDޘM�&��M��	�~nZq�dmI��K���MC�7TA&�8i�(�����GR�Zª�g�����h'r������c�~N��#�fw���;dEҶ]AJ�5p���'���d�:�Cώ*h��T�~��Տ �x��l���gRו�B���?)@T�����ၲ�"������"�.(�`���l��*�`^��Hh�5���IPn6P�4�)v�Tl�Sv�Z`i�Ǥ]b"b1�2ݬ��iw�؉.�1?g[����Ih����n��e���۾v�ſ��2⿓���(ߧ.�H���kbK���[cɃa�u�k��C��=�F�����z<F,I�!�9���i[���<7�S������>�����xX.��g:&��Ɖ�d<[?}�~��[x����O����O��tb�M	+<حMi�@,��L�$	3 ����o��.8�e-�ܦ�]ET�X?k`�P0�K�+�z(y���C��n�j�NPˉ,�M����%t���ߧ��PH�1!��}�-ߛ��l�IL�u�q��'���[�}L�s�=�U���n��V�X�}�^+cL�����r��ǟl�?�]�_!�_7K�c���*4C���֙�tݾ���J[���@�������=�<��L��7��o��;�s��*8�ܟ&Ͷ���J��Zq%�-?iꎿ�@`�}�}�2X��T��eN&#����y��wi�f�9��(t�BI~�N��@��_q��f3��i�&�^Y�z��a|{H�	ڤ�[�t�EC�ՀcB;M0�;X_��fbn_[��ua�B"4|a�p��B��\f��+&<c$��E�W~�t�>8��Q�S�_���ka��� ��]Pk���%��q!?���/��R��>���������.�]��I�Ϡ�]�m!���{��,:����n��]�1Ty��.��?�u��CnvS��/)������g��;�ߪ�WP�BE	��#���ʄ۹)M٫L/R0�uՈΡE)���
���)k�-�>�,?"�l�F��ˠ�z�	����.������5��$.`��'��;��2�.��}��Ѻ�"�HZ��!�e��x�-�y6��2�@��+iV����X-̶5�M�y�r���2����Z�Udtm	'�_��eĨ	��v�?_�CAz�>Xr߱+�|�#�տ�-��ξ0	�2�;�_�����lD��γ<(hCeJY�x��\N����)��Ҽ}��Ns����ș��㧮���3��Q(�&��pB�p3�����8++Bi��6, �s��s��Z�����Eӧ�Z�%��C�j�@}Ɂ�O�rc�ӺMl�%��x2�u��k��*̯��4��fM��m6+Sw��4�u��J=��'י���-��KH���3�gF \=�&f��?��5-�
l&$��!�y¶�KL�	����נc����Ym��
z�r-���3E�/��P�W�O�:��}�j������|�_BZg�: ��ٻ�U�����j�������'H�hҗr�.��
�k��l�c�y}�K)��G�!�$�� ���a�=����,���-�1E���+p��C����Ͻ���80=�qF�~,���hqu���g��\�M�9+�!�Ѷ�I۲�|���u��i:ݫ���Zq�g6�!M�P� E2����Ɨx�r�0lgf�.�#�<,g�qD�ق��42��� ����󩍜�Ԝ&���h�(W#��x�_*��k��@�ڃ��OW4�Q� q4W�wm}c�G��4�?�u�`,��)�/)�B{��41�x��$=h�`��(,9%���-%I����<V��D������ȬĹ$�O��1������.���8Z���~L�|��+ԺꄄZ��X9�>V! QmoO7.�'����9���4n?���-�@t�'���p�:�� -7r޵$�B�}�V?��Zm�G�L��
��x�m�|��qS	���"J��Ƒ�@@H�gd�tV45 ���>s���l�`��QbP���E�(��K܃
./��@��bA7r[9��=���<+����G���t���3�8�9��������A�����2Y�0�p8���1S)�J��{ܿ�5�Ѯc[\�ӦBZ?�y{�ޏL����]��C��g�>^[�ڂ�K��	�G�U��brn����N�>@�=?vN�T�+�_/!�����s�R$K@�2�rf��+"��1� J�V�A���.�߅��Ϯ�ƭ�F�g��b!p����(�mqcB��]���&�:i�W8���X/&�I�꒹��O��UJJ��Ц}hq�僑Op�1�"�+���5��"�hA�X���K�?������774Pp�_����w?�������4��.{=1��t'Bfb�Қ�pc&Q���&�LY�w7A��C��5��1���F�)I�`ͼtgH�V�4�&t\�{���fI����tH��+ �����sQ����Y0 ����m�QXл��~�fq���V�����
�P|��B$��`u]�6BF4{�� �D��Z`���&��>@p��9h�����oi��e���V�ݘ���﻽\ ��W�vǕ�Ĳ�`���l�A��e�5e��v] ���6謜�����I��@չ]|���}����
��Lʆ'��# ��˞?.���{��<��3IЅ�W*�%3ʄ�_���<U�^���8��g�h �Y�n�I0~zM��%�_�5���kW�%��Z6N��`�D(��5�������T�3Ir31��ob��J52`c�aP�	�hRYRa��$�`�lEּg3��I�^�yImb��=�o���RY ���R�S�S��~���<�=� H[�Ѳ�T��� w��8���0�1i�"d\�pqyM�ESk	+m@ j�X_�jY�2!����,�����v��� ��z5�-3����ܠD_���b9
Y1b��ߍ��~��ʲF�Gl�Ve�� @G�I_�W	��>+L����F�`�aB��Ի���͓�(^O��bR[�����7�r��'\���'�c=�9�\��<mm��u
���\��+2v�3�Y��K��f,�{�=�w��|��������ˇ�j����;���i�#>h�w����׿�5��k�w����9�C�kakC^gBFw� ��ғae��(l��$�ǅ i�;�$�W�:�IR/R`Y�X������L��]=}/^~
�WO�����?���dL���a�׿�<y�Ҁ��f�F���������Bg�q"�����I23Ln�����O�3�|XA���(5|��׆	?���~��ˉ9f&�a4
��}��9�=��Q��ǘ��j�i&jYh�b��2j26��hb�����OI3x�Ïd�٘z0 Ja4� KG�L����a4�%��	Lgc��-k3XԜ�-�I�i��+@�Lj�#j^�WYƕ ��[nx�d�p�2�E���>����{{OZ=5.�\d�㜙��0��b�xg�_���@a�B+m�P�^��s1��9��W_P|��7��@F�ec`�D���%�3�Q��
+��]9��	�!$��������կ~E���㌋f��K[��J������).����ϑ<��6F�	}���7��u������E"�NF4�1�	�Si�X����@U��Pr's��ڀ	��)=�y��~���<����oS��(�h(��d�q,bL�G�)iʴ�(;�Ed�1ߛRQ,��<���=�KG��a����8��9^�e�M������ڋ��}zwwG`��b�Z�������P�7��Mm��Ա,���pyy	�_��@���{���w,�����/�w��L�c�V�'O�@�t�8�9����ue�Z�������я?�H�S6O3�V�a?c��yj6&�|��a���?��5�Ѽ�ɥS����F��]]S���ͷ��fi��%��[����H��'/ዯ���������z2���g:��`�D����=j-+x��x����E[gF0ͮ^��O���O���޿�lnJ�6Z׆T2�X��0Z<��͉���*����h�Z�6�D"�s�IZ���DX��P�|�ŗ�̾��oD 3+V���$��hH����?����2�Z�U7N0�'`���|�T��5t�撤�a#�%���95Lzb��d2#M(��e�4LE���5��V�}�p�eN�3�y��0�
��_FR�p�ǐF��p7 j�וࡩ��˲E����DpJ���t}�b} �l�]-����ZD�f�t+�X	��ˊ,A
d�(@���|Qk�`������uR�1y���$�~ٌ҆�
H�X,(��=�&P{k�����aMp5��~@*�\@M+�F�¾(Yk��\�&���w����}(nm�I;o*L����#�HJ���9������\��i�k�~i�B6z`���A�ޓ% ��l۹J���I��S�;�y�J0��w�{Ji��McY��5� ��<�n޽'!s���F�}��+ �C0���f]H��U�g:�cC��
eY�^���f���u����m�+���yL~���WW�0J��W�n� �_�y����[ �- �~�)�$/`26�$���/>3|�(_�{����|>=�F9"��Ɖ�d6Z��5q2|�pk&�aFpޘ���?K�Jz�i�{:1���o���va���9uI��Ȝ����~mN�[41��h���>��b]Ȳ��-iXȀ�����}�:�8'�Q(ppVV�����b��G��`L		ׄ���I7��� W��w^=���6�]���%1G�08J/�H["K�i�9���nQ��^�X�][���G!�*���%��h�F�Gn��2�=�p����;zg*��	"�}� �~���!�	�u��]�*�>a�.qč�l|W��l"���ɪy�C�fl���:�+I4j��6�@R�x�7��I��rP���ޏ#a�^S��[��ָ��H��:��/K���a��.��*�큀����j��82eiW}�lyI�{�4@�u��r�o����8�q��%
-,h�O��5ƫ;��ر�-�Jc"�㣒�Ti=���M+�����>IB�M������ܶ��g�s��Xa�2�[�B�D��pn�;�4ݗXA�������]�+3wйg^NJ�)t��Eĉ���Q�՗�����`�Qi�:��t'B��o�"3/V�葙�eSp���i�k��6B"ɑ)R�œ��:Wd�%a��b�%�~f�����sojf&)SV�[�	'���u���?ܼ�z�2�;D��Lja��N1���I6X͙?5YU�J$i�J(�-�ez���4�̍�'�ͮe}��91���F����h��kx���f&�+)�ؗw�,8�o46��� �ظ�͚�U�Ni
MJ~.�s׫|���w��.�&�@;a��~5��Ob�v+����ˊ&�|�}�eC�0J��v���U��(XK
�q�d�t���
Ժ�.��"V$)�Uъ�a!�� ?�^?��z�+WЕm�&}'}/��on,
�AbRR���h(����F���u3fK�jc�o���	�R�g��$f�w-=F������O0~�O�<�QH*UY�4���{��PX	�S�MY�A��y�i�/i,fxW��X +���*$ �����v~/�X��9nl<��6�&6Ą\�nL5����):�B�.���ň���⟛�Ρ�y�8��ӝ�7����C5-��~��Cn�b�ߟ�(G�3�8ZmV	�׵b_}�+��#~o&����S���B�W�T�o��tQ���(àS
hD�al)f���B4\�a�+���%V�d��nO:X�B�k�~���=ECs�"��ܥ���Z�����kY�ʜPd'1C-��jSY+jF�;��sBZ%Ԋ1���F�Eѯ�5���fwŋ�3�[�L�,�޾�L����-��.5gLȿ��$r��rR��*ݬ�@a���h�)����#�t�ab�!��mk�:pB����?pW��AEK�v?5��$����ll0e�/��n�2�ú#�N�(����;������f(7�����3���fc��Dl�HS�u"��<J��q!���������BP�BZV/��n��-V[���	JV����~�� ��c�$K��f�W���<�y��`kb	v\R�7/��fƚ1�*]g��Jy�G�,Q�+͑�3�" ��k�fɸΟC�x+�*^��ݒ�׮n�n
�K���'���h�1�\ �mj��s���D\��KQed�C�OA ���k��1+Y��*�Z(�s
6�/�̤��$��7�vG�[c���>G��b�8�1*b�7�l �]��,���J�#�l����ۧ7��F�ab�ӷ�����LD
���B��S���V�LHH�R����&z ���l  	��VHs�8�ȐTU��i�K�kձ�f�3�Q֘�C�l��B��$	�����O�����X�Z�,���'�`P�hQ�`4O��E!�Xk�1��p�� �����y*���)���хzܐF?��%�f��ځ��V$l�_O�et���g�Ej�vY9�ofoɷf����_$`�M���5�S<���U0 ��]]"�D���|�ɤ�C3�:И��KJ]K�|��_)׊r�H;P�+�M8�j�ܦ��g�����c�p��\�(����Iq�I��@ai3��m�\B�2���-��5�@*K�- j�6		UT9��3W jk�����s=��f�����pRVn�a������`n��]�-��϶���Z� `E�
�kVA�&h����
xS�����
-����k�!K��oA^�����xg��R,�F�Q��/>�>��g���?�G5βM�p��8&��ƉP�fS2'9Y�A-��:1����	��(�_M57'��ׄ�����_Yi�I@S�B����6#-]-9(���1��t�Q��������>6��M��Ċ�8�vp�K�o����������JvE^f��#�^Č��� cBsv.�)g5��F\�����j	�,y#�T�(��ɘ5�`<b�Z8��B(Gk��oZ�a�$����*�����t?-�lX�Hł��6��O��u1���Fʬqid	'Rw��׵r�q���߯��y
l���q7�6���f��V�:~���xq�(�$�@�I&�Y�% 8�H�e+k*�|x�5Ժ���E��LFȂ9�Y(A����@�`3��\���n�|�^��Ь�:e��f�5��� ���!��ͺV:�
(V	�%��]&b�#���a��R 5�{q�ʎsTl�[��kP��xz�L�0�bhk9���T���ZQ�`�}̟
Z)�[�U�q�9BO �c����e�~�)������w�8��'ɻ��L�l��4�ŵ�s���»����L���	Z�r��ɘ+�?Mx���Z�B�w�&�b�܂~���9� Di�A6�����W�4�����x	]2e8���)@4+р�==B�BʐO�Z*��i�vp�6�'n>q b������9B j��p�	-Q�i�+1O�9�c��*ZЏ��c�=�q��9P9�/�v�9�FkH���U���\���oHߡ�A�����A��i+��7�j3�RY���.1��w�ؠ�P�:�?yB{5�6�w*+_���?D���˵���B@F�e�n��ZE��q'�@���X
�� �|UB���i������+k%�`�����������G���X1�����O�WZף�V��"V����l`�6I�����e9�`���h�B�w�.�E��lʖ��i:&�N�ɔI+Z��DyMv�b	)E_Xw/'tC�4I��}�̭�9��c�0�Q�غ�1\��*L5��Q`~G��߿���j�r��h�7� �#�l��7�t��u3oh�E�J��VҚ4kiR�Ot��I�@��t�*�F����	�^7�~4+k�5ڐtҬ��4W�ZT��&���@�v�h�\s�\�$̫�@��+�Y�qrF�zkz�Ѵ��洉��8➂�Tj�DUͰ6���d!&IE�d���U�!�x��j���P�~\>+�(�?�+LA�wV�����d�v����+�]�Z20�����f���Y����0�w%�-��.��0`;��n��|��b�/�maWY����Ǧ\�X��c��"}S�n���3� Q�-8`�N�ⴶ���J��ŰY;٫���V�"(�MA����֕������+�C����m�^����l8�`-�4M1����c4�M��3D�O��W��s�$(4�u8��c��%[+�@a-l)�A1 �|��Q���C����bsg�8Z��\�2c��Z^�2t�tGm�qC4�ѽ���̣?�����Ï���0ɯ(٘QZ������3Y:
�8����������a&�������,`�N���8��d�L9�e!YS�5s��^4��Z.(M�jg۔�a�5�"q8�u�Фg���T� �5V�{���CGN; ��+�6嫭;���v�*۾D������75NH����<Y�=Tf�E6���eO������x���.fu�7LF���oIrW����Ǌ�>�_f�_;��q���� ���k��B��P;)��b|U�XK(����en������2p6���q�kO�{w��<��(����J�����X+Ԋ�����Zk(�uD�,��B�6X%gxM��`*��X�Z+i��Ի�$*�L^142|�ͫ�����z�+���@�Wp��b��6�}z8}���_|g�4�XE�¾¨|\�f"��V��1b� gт*-�yx�LAUvUn1Ijn�S�Tv��l��&^t�/�����e�A�uM�k�y����xŒ�@���}D�"�ڕ��A��D�c�  ��I�<F���Y;ʷ�'$|�(&xB�o�Ba�����^6�bT� ��'�s�����+����~�z���N�R�g�@���J�7��+�� ����qx���zP8���I�%Pk��J�o'���W,Ѫ!p�o�������n��^���
7��Z����`�킪^�Z���XZ�j��2l�W���V`]���)m5M���
/��2�xG��4_n�B_Պ���R�3��
�Ù�Hg7ʉ��FS�x6�,z�O ��j�t�4!���NH�OK��@�Ċ�$2�kiBW�L*�M�9YL��&`�A�H��L.	s1_��4�.Sn��m�<�j۞��Eu������A� �GeW����X�u�	��RyOH:+��/��aM;���Z*X㋎������-�	$�Ų*T�8��ݧ�D���b�a+׽�ӵ�@�R�M���-����|����z�ߚ�cj[�c�%�*+	��}m�!�]�jU"x/&kU�lb7���Dq,hN�����V�sl%�]'��.��b��K)
��%�p����w}���3��`�d���Y��ٔ��߻��r~��Ʃ�I6��� �i��ت�7)#-F7i�+h$5s'��>��T�iX	 Ѽ��j�!V��)�iǎu��c�h�nb��-@G�f��7Ś��>�M[Es�6��b<^nl�IZ�qu=������*8T��ePp���k��.�)�j[(S����+Pb���uЪ��ni�����ע�31�V�)�������SΧfw��غ���*]�a74�@���o[�,����c�k�$��ߕm�^����-�8F�]��A����#�Q2�p��h�<�Y�U����^�ul%�%��.��P�
�d'��gm ����-����߾��b�������x<���Bg�q:h �I��V��50@��O^��/.����=2il@��� ��Z�!��Tt�4�=���s��K���n�5'��!
iLr|(��G5U߂���ݳ��թ���Y����l�˖@�[����c��1�Ϗ���.������ͽ�}u;v�,��ǅ�;�>�xE��+Ide������SYK$��J���9\wE���v�z�B�4A�W����wR����U�Z	�ڣ%�_j�Jj�r�x�-�������]��XA�
'l&�\�ᗿ�%��?����[������wKȿz��FO�D�Hg�q"d��
�w��nx���q	�Up	����A�ߜM��8���|̺I|����m2+��mF+�E���a�I�Z��A&vf����d�."k1n^���P� ���y�\�@\XԈx�
����.E�s�]��9Nu=&���:pث��~�<���ic�y�!�����k�~�����%7�@�}$�ɵ6�1Q��S\�m�o����l�r�׀�Ƃ SIۅ�4���8�X�Z�Jo�-́��#T��c=�es{9���D�҉]=$�P6��@\��>T�Ki��W�8�@[�Ru�r\���_�-����������=U�e9x�i ��Ɖ���ի�d�ws��G�E�ޔ9e=�1����p��$7�X3I�Q6h_��K3F[9BE�Y�q����۔��z�1�դ�F&_�9�̉���綆9��bd��R��[�&��
�Vy��=<�~^G}B�v��˪�X"�vm�������u}`��$&"vn��m��ƻ�{�n[���ϐ�Ɩ+)W�9�f+ވ>9�����j��E A�Tm�p?E�'�"�� ����׍[�>�-$��mk	�GQj������6T���������[ ��N�?�{Jh�0�o>�,���te>W��/hW���l��b~\3�#Q�O�Nl��~.�����Ϋ2�o��S���������q%��.��JD����N�\a�
�������� e�K(����i;꥘`�gj���^$~�H��f=�r��ZG׏�t5�ڄ
��%n��3��\e)Y_�b�Zꢵj��p���5���0'H�;6�,%�dih�`A9P��7궁�ݱ^��P�*>#�I���5.�Um��[�d��Pͽۖ/���+@`an�r~�X
�> ײ���e�/�#�5��r���X�@�<������}3�0Y&G�NǼE�䪑���l
q�:R-eA�M��1JN�������4m���O��e4������xki�J1Lhed���$b��l���`x�,�k�I))�:!aGº���c��X[�*!T���$�%�=����5��1Zab�
F�Di�I�g@?Qw2`��s�}���)���7b�o��������A�b�Z�xGI4��h�W�IT۵�Z9�EY��`Sg:ʗe5�M�Q����M�.fyc5/�gm5�ا��}ӯ�,`�� �v���A���]4�F��~�-�Ш��ois2/v[��mkM�`�5þg���'V�X4ܝ����s�
����?��BcN�vH�i��C�o��rW�{�q(��u�j��X������P@���-��>๊R�s|Xe���tfY_*�X/�V�0Z319��T��VV��LT6����dj�{I+��F�QOǜ��ay��J��p���ɀ��v������`��/�����5|����?�&�;��O`C���6;'�*��k_[e����"%�����%{�q�����ܯ�u��޺o�z�����vGW:oaEe�M#����M>����� Va�3ѺƳ�H��K�E@C��h��s1~���g9�S ��:��б�/�J�ra\�1[u^@B�U�����wS5��D��XM�~Ӛ����t��QY^�ls)�^�eA�� LK�19nQ�r��e�
��%�7sZ�ʛN�.���41�1��}�{�T�*?G�I�e�)ş=��F'5����*7n�6�L���'���Sx��%,W��BF��H����Yq&�-�dA���U�sBAV�f��DJ<dܔ5�ĕ�n��v�Z9��h��a�B\sR6pS��[h��5��\�-�c��}V�Z��4O��3ǻ.��W{��RȪ�_�[L�*����t����u9�}CbC>F���2�>}J���F��A���*;ֆ�}m��\x,��ڣ�TYs)��e �-�+j&*$4x���7qDVgseHn����9@��#����w�4`���	8��ݢ� Z�� wa�)q�-��h��i6��:�F9"��F'}<����X,���~~��R�U�B_�%�i	y��_�����6��F)�J����H0��@�"����h�DԳ�CV�$�~�m��7��X}B���V�[^U[C�ͼ��6�����������~�}���]�,v�[����9!��SG����\�[t<%�h }���h�$����C}-o��`X
��M��ӳE�GZ��ƛ�� %�2�?�1}��NIT���6EdPBAڴ[��m~g�
##7I�r���pI8t��f����c����f%�Q��R\�gX�)G��>�-�?���6�Hg�q"�������u��Û7o�׿}�$�����n( ��a�ź�@�ژ786s0�E)�WŻ�j�W֚m�F�^�R3&'p���֙��w3bQS�Y(�xv&��^q��߲h��;������.�68��sǸ�~��C���]_����߭��_,����h/��oߒ�ݨ�[jIq��Y�e%�c����{2�$+F	+/hŬH]ɨ��΀��*'��|E�M�mB��&(��&}�+�L�W�8���n�h%�����f;ƽ�F�����/)`<�0�݆��>�4�tnέ�q>��LG�3�82��a:�H�
��35����'Ӕ:"w�0jW��̗�ٌ�F"s�z�Af�t*B*I9ۧ��$�[VD$�Iq�5=v�X��2�q�l��u�G�	\f"�L���=4d����	�r��N|��1�.�j�.V��{o@���]�l����G`�����=E:��B����
>|�@���@�!�u#�/��� �  �n%�
��H\4����:x��bk��-�i�B�65��yxP�F�n_m��5Y%�Z�S���o�	�T�M��\c�@+��Y�(fx*nh��
���p�������3
]���ʄ�t>ӑ�6N�~��_��u���g�}FL�W~�I��yS6�+Nţ�EѶ�9�#��qY�����4�u&Q�D��v�ʮ��m�$Y)���IP�k��`5�����b|���瘏����=����R��\!�E�=��[N�`�c��2]�'�u?��ߵ����^��W��h�����!�V��WA�o���s�O[6��I�����W���v����4�=�q�E�V�T�P�v����<��E���֏JC+Gc�h���|���p�_�Fjxge�FE;�b�D��A�0�������'py���xY�,��8�Q�Hg�q"�ۯ��7��5��?�M�,OI�O�py����M
�Պ4���J��cւ0�fŉK
�.l�� +@��7����	�U�b?؜���,$��49�1	�&yu�������`�?4~j6�6��$��0%��֥�m�-8�S�uiP�\K�i���]N�+m�̄��7�L>sFf��~��Q�[y)��������Ƚ�/֣ϝ#��e�ʌYo���֮���֧����q���c� ��Y�������V4>��>���(%���U��Rze��=�s��-%!��$��k���4^I���JA�ή��ǃ�Z.��`���"���	^I��-���\�a�?D	j"P�q�����LQ�(*[e�!��$��%���QV���9���Ih!F�{sWS�'�O�Lǣ3�8z����|>���� ���s�ݢ�9�#�R�g���X2�6P�	�7+D��!���=y���'m	/I�Z��<͒�0S6k[(F�B^U��5����٥g�4�q���܄=�M����hH�J�i��5�zۤ��~�����o�� �~�ې���+�$�3��jv5��u���8�T�C�=�� ӡ�W~_]wi��>i,/P/u�1�Z]`+{���X)�-G F(���)gW�J%�9�x�����1�k�0�[�m�W��X.j��x��[�j(���y��z^��A�ALe�Q��ޭ�epo�����3O���t4:������O^�z��K�"KF��N�E���Ѱ+�/�t劄=��8�0��Wͭ���dӧF�a�	2�F+b�V���	��Uٍ�J�PH/�v��Vc3�Y�\���Bj�2�O�JTs�d��TU��C��������n�d��d$�S�pj�JW��i��<@b�C���9�%-{W��}4�j��s�4L�b��Q���	�n�x�{��Ы[h�4��c�$<Ʒ�I"��qN��#�!�(�JMQV�ƪ��}Kl�'Z6Ҝ�6 ����E����?�����%6y_Cd�@�F�~*Gcz���(c:�߭KF�6&̦��rcÏ0�0����9\�
=�~D.t'B�ʟ�U�/�>�5�Kp�/�6�-H$�uf'���1Yf�KS#,�����?Q�Lb���[K΋Ģ�1zڪ��5����N(��c�a>1H�R��Oܩ���뛝m��x�i�KJ���1šb�nO���b�3M;�uwݮ�.7���j�����;j���*���. ��������k��Ci��~ȵ-�U�{K�[zr�k�����B��v����ߏ�}}��Eu�����)VB~�I�*�#280�r]X��  w��XJ[JT�ֱ!	����؀��b�dwXi#�_�����|�$��r���H��F����ܙ'B�M��^ ��+x���\���+�6d�k|�9Y*��%B;��ƕR�]�|��B�Tb!��K�f`4�Jr�<$���(������%�I���MON�1P�^�և�-��lA!��m�(�M���h�Q�{t�JB�+�Q��FT�#�գ���I����i����н�񡂻��c�>n�]�֩S�:vu�� C�������Z�ض�l[�\��>h�{�3��<稌JYjo��E1�X�ĮDQ6���������n*l$���ϣ�
�e�Ȫ�g��FR�*��P,%��	��{�<}��E	�ɢZ��p���l��~����e��
�\^��tb�lIe�0�?
]r��2XD���hvTvV!0�l�B�1��ʺ�G�$袵�1���2L"K'���./k�$���$��p��?�� �ޕ�ّ��]�������@�,1��b��2��ae�VX b��իg���4���M7�}M?���4D�"�%����.�B_�@��?C�>&�,K&c׻��Y�b�`�3 �F�0~�R�!V���U���B�{���Z���M;�\v�2dݬ22ǵ�o?B'�A%���9ם6R� >��%4����̛w���ج���2�dS�Z9ɼz����ht'B�4-�Y��������ۿ�����2W� ��u
ݎa�f��@a�
إ�ls�-�yw،���1��J9����e��C�&ʤ1+�5��� �;���Oܘ���֚Aq!T�}�>J�v�?L^F.�V�.awm�M�e���@,�PxY�ę�yZc^�1���`��2��m�v�6vW��q����D,p�G�b�	��B�w���AZ2�������[�h���{<�-���k��U^��vq%�F�s�z��9`�vҒ��S�2T�ZMi��&&��hO�=�A쒔Pxdic?Jk=���	�N FK��c�LkG)�.GdݠyZ���8/}="��Ɖ�tvu��Z����Y777���p#5Z�Q����7��,�����<����]U]lv��&C��Y���I��8� ŉāF�@!��Ob[��$0q,� K�5Z'�%qh6�=���;g�^k���^�*vKE���x�^������^{mIu�dR�b-���fM�,�Qz8�*���1��#�� {n����x��
Yp�A�Zɮ�E	�x�D�B�sFx�EL��.�Bo�43�a�S4�Ǔg$n��^{F���qI�¥X�4����OŸ`V���2��XFa��o�=)�rޢ�z^����G��r�Y}��H�H������&�A����������?<鼖Ϣ<�����o�#g#.��͘�g�(�1\��8���F����Ϝ���]�F<yo΋���Y�~0n����n���v)��[��b����\��-ܭLe�le
�,��l*���� ��l�"��e37+1���j�C��u:xQX��kdɅ}|����|F� ������n����LFc
�T�u�"��Q���T�x5���"D�oZ��`&x�Y����yN�<4w�	\��`�7�g'�Ń�T�{��{��WT�P���E�άgw���zx��W�t�fķE�ˍ�峤V\	k��44�������)@���<�J�e��*جb&%��=3� Qs�<xz��P%� b
w!sV� ��c<v����BiȂ�c�b�bɫ�";�{\�ԙ�f������F��(�"�b�VϢ4~�}{E�鴁>R_����E������I۷災�"?�����}�3���2�v�{S�E�^p|�$pʩ�t��J�sy�X�q�9�OY�DΜ��b��)�n�8D����46 ��~^^����io�Ɓ�'��p�ka�g˨���\�)�u�b�Ԫ2���tj���y	4|�M�tZ���	�X�2󌸙�$]8�e�hn+r���҄�@���C��>�A�#����JN��X��+��>ؗ=�A��F=���E��S�.��3�a8K����|74&����b�	�uhE.KZ�cdb�Vc����+5V�,��sIbDNޤs�l�53�v���$��_Ű�1��\'Yz�S(E�r�n�=K�H�!O�(�7�.���+mB.54�'PRL��!���*;"�p���kr%���г�]Ԥ�����G�����Qy�t��;��R@.�S�+tE�?���3�Rv��7��� z�q%~�����\��5<�3�<���%B��\����y��I���.�p���jā�vƿ ��}۽�,�\=�矎\�wh,�\e��4�*��f�c�� 4SŒnэ�������%��N����9w)ۙ�G�㉮?�ܥ2��Mf���px�,��{��z�D����;��y������7���L��,�u�Q�����(�J�D������g��$���D.���]��gdSϴ1��e2�%:<5Tu*j2����AU���x橄e���G��O�靥j������ ��F��	L=/cvF�q�^�)��_?7Ia������V6fZ.�x%�J#��ZW?W�A��*[|C�o����P�ci/�*t�hd�<�4q�֮�T�p��p�ya��i4��U5Q߅�m�[�-B�~E�\�	�'��E���Y.��)�<�U/������{�%z�^����q�����9�sv]˿=�,��H5\<��[�+�d�����>�`���JUHq���1K��Az;�����3z0��ق��-�_	BDJ��a:�dqi�˙c���E�4ѵ�H�R	+��De4��g�����!�b�Õ��
�?��Zyf�Ȋwj��Ѧ�}d$Q�::�2FH|.CY�3��BY����y�X�Q���Ɔt��r��%ypp���*u���4���lE���D�ñ
aU
�ac�|L#k��>�K;}�[z�e�1˓
��+?C��\��>X��LL�<-l�42�E�= �\�8���ox�ͽ�V)���g��_."� Z�gs�r
̸W��2�k�]�d����[���7r��г[��{�xW�쫞�#я�p���5 �D�a��NV��KM?X��<���[q�p}��F4N�'��IFy���>s�9�ߏpΤU�����9/m�ʧ)�m��[>��s&F7w�H/��Au���j���)�g?yy�'�e*�$js?������.���lƖ�l%��(���e��d,ع����g!���+5�j+q](i�觛υE9��<L?@�4)���$i^��Sqs��)+}f����Q����w�^��z���)n`��t������\�<�=�� 
N<�g���̟�d#_*�(�MH�,��.sE�3F�ݨT#�4��uR�x���إ(`�{:B�I��4<��ܒo�	�g����Ֆ)
��V>X�z�,u��l~Y-RR�
BH��iCQ.����Z,>�Q�낯��^���
y�h�]\���"��̯H�#&�&O��aѧ�3Ie�o���K
�Sa{�[�~e[���?H��qۣ)��۷XO:O���~Ǎ{߄�8v}{6y�;��|�=oe�E�^���Y���脜6��qZ�Z^����L��n<�DC�x��u�Rj���=M�[P���
�WJ�S:�ڜ�S�xF�a!�`�+~b1B[O�r� P��4DX�}����1Y�:�ayf���_�Z�ӄS�0�=Fy+�w�ެI�Y���9�����c�)�<͒4{�H�b���wl��g���_���͛'�
[�W+R�5H����(!�4)$��o~IYN��H]�4@"�D�$)�=Q�S�NU�{$A%)�G�L�z֨�r���$��F!�[�3a`$@��=�-�\HW��z�V�WK)qy���pXځ�=%Ν�9C�.bQ���	�\������yn��`P!��>n��{y��gۙH��2|���7���^���}����3�2�?��,p���b8-z�L�<.��H���q��qQ��b����s�5�ϯ��~���sf��`G >̓Β�X��Y�y�H�&;������~L���l�\W~{��s+�~�-A S.O+���^m�f����,�>�l�t�Ҋt�(�UF"}r���,�{,���` ��[�|�E��ee��:&���|/|}�CF5��T0=G��Bg�)n��q4���������[�P�+B-H,Ș�F:Q3� �{���
�Ӭ�0JF�ЉcR#'��%�U���4A<��2Md4��:�<�5I�+�W"�=8��Ƙ��S�;.C�^��Ȟ����Hr
�\l,ל�W%e$�-$b�Ţ$.㕊����8�{��_)׽b5\�8�Y����^�.��xg��td�~���G` ��n*���$uy<,�z�$+R/s]{��L΂7N�gg�cZ|��Y����.�+������)��<��;�Ϗ�|g�ǥMhD�Y�w�$e��*/��2�b(M�:�"Ήt���l*�0��|���{x΋�G��w���n�g^�3Z `�%��e�C�ts�2�b��}�iW�@h�99Y9;�7~�Ȧ.���[���U���xVE)��[
�-�����jl���_�3c��㟉:-�]���8�9~�U�Q�U�$����-�'4ak6u�V�
<Rϛ�i���]�Q����h�q(��D�s]��n�F"��SF2��9�U��)IZ'T߼
��Zd�֬K�Q��d�C�fKZ��D��x''��XuG�
á~X!I�+B�#��3����{�.����(�3���o�ɑ$�'�jƅ\s'����uJ�T�Q1�[��R���Ȟ%�y���w=\eB܁k@g5�%�t����f']<�n���z=������b}�0P)�|��&q%�d���
4j���'������C�������3��=��灁��?o��qQ�;�"-u�9x���Q�p)4���g�j�<�d6MX��*/bS�ۈ6Vc�{�2��.�W�%��k�(N��JD�ܔN��Kx���9
����Ga`4�V�.��-��J���V���t(�z,y/�x[e�����=�,���~�D6d��焿L5�3 ��T�<~<?	���E�wu�X�I[� 2pD�E�D��T��6p?Հ�F:�c��V,���.��3�����d>��X�՜D8b	⚂���hB$A�����}���� Ur�-v&q��HE�^Y�)�'��Ԁ�%�L�I"q5�"H�ۏ�Q�ys��W �7�#5�V��(�+�B�,��+�ǵ�o��}�*u	=.��8���u� �aQO3aJ��J����Z,^.��}��<X��L)�=�&�L��	[� A@�%6���|+�8���x�{N?#@c���ә�,��6\�rQm���3rވhdY.�\F7<�Wƭ�g8���lg�e��B��w��^ؗ���q_�w�̏ٯ���,�v�R��"ѽJ�|�v��ˈQ��R�{U������܅E�(KGO����)�}�a�� �gu�1�8�@�s	[� +�aՎ�s5�z׈Z"uVZE?�R���R�kI�2���#��i;��)�f�y��+i��y�ѫGZ1�LЪ���g��l�X�+��c�:�u{fE���ݝ;�#D�-�љ���X���5�u}�b3�~�/����X�k���i��Eݏ�Ұ~d\�����_�f�� ��u��*����Rכ,M�����Զ��l�E�~�K�z�!���ZCuEDc>��].��.�fS�|m"�.��I��Q�'���D��N����d>�	��D�(kPh7�:��$X�3J�W�Ŵ�;��̐h������X�y
�<�G�*J/��R�bL����\a]`���/ĉ�/�7<xY~T! BЕ�=9�Qq�����B���CgaS�qY�-tKBߪw,G���@m
��A2�Zn
�Ł$��(�/��\�:��R#��Q���4�J٤
��ټd�ba��������.�����ҼEߌ|Uձ��<���Y��
>���v�~φ�O����;�v�y�nO��3�u^db�K��v^��U�eD��}�*+�3Q;�ϖ
�ԓ��
'��<�3Ƙ���c�f3+'�����he6��2u޼(����>Qc�2�j��:�kqŴhr˲�C���Y��ƔozLm���:��X��AG�
�N���qbZ�q�,�&N(�,�5���2`QP٘`��c8bd@e�95":0�kp�݈"�l���$A��*d6�2���V�VD��*I�w蚩9��(V*y|�������QZ����i���A�)n`�����t�O��N�{L4�n��G�8��\��9��x���S��,*U����ck�W���}�ALO E�����K��A�"�t�g��c�������H��T���(��7�2��9ÉE��y权Bé��ҧ��Ft&%pVv �!�Ff�>=.�k &Rd�#>݆;`mbA"fH�b�RX�J�l��>���Z�DQ�"�)	|�ʏ�J�ι�%9ȃ��h�\�Ƣ�(��P|FK������楨�2]��{R��bs	������ᬑ~/���푔�
c5���i��x��1V�"gI��G��~w�A��S�}�}[��}���I��H-��s�!���~6�,�WS�1N�R�2k%���U(S3��T�zK�'��Q��AT",]
eO8?��1��9]	q"_9)�giY�q�gb�qV=FV
�)	u��(Ll���_�,1�bGE��*N2\CC��&�s�����b%�X1��~B�?�����yFg��	C@�	��t]+<��*��fmQJ^pw�L���q��\�(_�~��G�k�"��:V0_)��0�.���]��g`KFq8�7���eE��1lԪ��u2U����H���Iţ2���.��g�,�<a�#±��u2!"��#�.x�0$�)ԫ�Ø�~����2E����e�b6�
&�.���gBe�k�$��"����Ђ�� ���0�v�z�g���fM���z~�� 4EB�W�� ���+���� �`�0�ff�U'��^+��Y�:���7�*\�\��X�-\K��H��?#�.JyF=v�^
���H��R�q������?�� f�޲�A��E^BrA|?wFhiP}�8-�V�g8g���z��.���EDV_{\j�qѐ��ܹ>��w}�۲��tڇ)� X�79�z��+�>}�ĥE���HP�ץ^t��z$�vPgB�CZ�Ǹ��!U� �J��o�ʬ�ӹ� �R�UUY����̇.��5��غ1�k�A��Z8�����g>�D�^e)a�vy�/��t
{BzV�Ͷ��0�k�}H�d�tL���q�'�� ����닂9�`nB����0�N�x>M�"�&1B��F�g�Lts�3�9�u|Ώ�*87�1�#t)T��z��2ҥ{��[9�4�~�h���Զ��lQc���ރ!�D���{���H&C]��D,�P��T�� �0��d:QG�`D�#k�6N�H'�h4�AlV[�I��MO�V��E .�4l���"���h�����_���t2�9T"�h��(���cep�uF(,URxsF:��@Z��^5��y&诀�r:���<ɩ|��Y)�a�EA��
��j�T��S��2.���.��yNe�[�/�/#*Q�$��;�󮬤- ׎�$�.R1z�&�%��,;x�{3��Ӥ����Ca)/1i���ʕU���J�Xz�N�9\ڧ(�����M[�i��%w�ԱW�g#g�22a�����3�%��x$�q�ﳽYΞK�)��P���4,I"�vi%RS6+s�߅�D��?��wR�#a�'���kM�Bf�K�P�	�ĸ�Yx�,-�1�1����_H�"��Q�&#�	Q?�_�g��L]y-�Ƶ��c�i�_�-z��)��(���f�D�r�B#���Az� ��yN�����׺�F��l�E�2��ˢw\�iٖާ��P���jň�z���2b��O�p�t�^��U�aʌ�S	��r�<��=�o�c���x�>�����.|'�`l<��l<�z��W+o��Ke<���qO���2��t2%���8����8fň
����JT�	qq�'>��Wk5�ިKMW���S ����ـ��mf�1�f���)��wpp >d�4t���|"z���q^Q��v�C���)9�� $�E��":�L�n�#�b! ���H�d4WG*x-z���L(���t�3�DR��$��@,�n͢��'��r��j�U.��,!6�s8K�*6,�H�`��d憮FPю�jYF ǀH}P]�s��w&�(+��q]5�Hi@	����Ǭ��})ΦV����]����xR#6ʬ���@��1����sW�,"gqʓ��lJ��� `++V�g�� ����`�ݷ�*	W���؁N�����y�a�>DlY��R�3��*z�xK-賋ku�tnv��N������A��
���a9W<�˦�[��������,��]!��^.,I��q��l*�r��h��,D�x��"�҈��Ԋ�|���e��P���,��,�;�y�u�UJ	�ttm�gZA��?��ui��Gd�l�s'b�)�������p�2�ֹ�ay]�o���U� p�=��\�9!�@���|�Ѩ��FlŅ��c���lG�C�׳z�*�f(�[]�y�#�?�Qy��O�p�(��K�=<>�Z�a��� ��͌LWkl����p@���ֶt�m�\�2:�L��IG_����;:���;9"����y��w�5����\���G��W�ڵ+��^�-ԧw��\H������2�����FP���ܻ�����,�6P�R�k@)Z���b�ei𒰿�{�;��h�WP֗�~g��
ׇ�3��G��3,�H�T�5�zVe�ϕ1�|I�c0��E���?��af�fL��:��@��Ȁi�}4]58��}R]��+�E���ƶ0��iށ�(�-��V�,{g>{VO�t��y�#���h�FqM�No�H���I�����
8:(�����7)�2�^V����r��Z"��T���8�	A'������/#T��U"{�c�WY�W0?�g�aY�4�|Z0u��""y�3��y�eQ��?7�q4��y<�n�خ����c�η�>R�[F`J��{�9��@�y����(h�!K�I�;�M�?�0ȳ��c�zh�J�b"^c��:�5i�oa�P�F=�y����aHm������&���-��>�Y��kH�^gc���;�s��Y���	���?�뵄��Y�vw�i���Ha�����6���B��fC��U��I�
l����}�����u�@����x��`'�ڞ���9���p �t�y��\֟܉i꼧��p�*x6FJL��aRݰb�(�;��Z#���9
��3�,B�:�Ӊ�"��A&�x:�Ʋ�wWQGn���r��|�����t�+�8�2��:���#L^T�$��,Z�@~Qc�{V���w4�HW��pN�$\�h<�v���Mu!��g2���tQ�Z�k�.*�i��79)���Lw ��I��Y]-l���\�p| (A�C��Ш��Z\P�]���Z-~�w2`t��t̓)�O������Q�'o|����;������\R�� �k|��E��-���$6�TIf�#�rW�gvof)_,&��JNa/[oKm�~ZI#��-;͖�浓��\��إl`��\V|���� �+颒柹��K�5:�|+C���}�[�4�	�І������(8��~1,Nq^��f9ŮХ8sQ"�WN��Ü�����,eF4\�(VC^��0���"�;W�����ݽ_��z�H��Th s5�hG����l�dmc���{l +�8&�m����V�ful�\�j͞?��Ї} ta���}+��9�<�Υ���M���9::�3�>Kp������l. ��R_�$��³A�����y�uh6)���o�:2�p~�� �jE]�U(�n�Ѵ(�':?:��^o�s�Ç������E�
��D�u��Wc����klp��3kk\g���Ç�mln��v��1�u����͗�=Щ�䄉N��8<��l<�/H��w����2��_��N�u5Dj���u18� �b�˝;�$�S��57uA�Te�]�j��֬��z�X89᷶�4lH�����C��{�c!@8�Zor�<�?�s�������G>�}�&:����N�D���K)^B�H`�j�,갷w��~c*��^�g����;[X�m�J`���z���iX��j��iZ����<Fv���3^�v����}X�@g��:ñj�꺀���a2���N�
���G��Ғ�K��lJ:�0���.��V�}Yz+�&⥑��d3��*
�
�^�d&S��s#ҁ�ϻEB�'../�N�ff4>�f�>��z� ��Q�:���������֛�rA=FU����w\p@�b���, �JI�,�.�f�R"�g�mNc��H�އ�gB�rn2��`8C�?}D���PE��~�r?�9x.������5-ϕ���G�^���T��#�0�I^ľP���4E�tE��Q
/���S�9y����'Cv_�޾�c}��V����*2Q��Ѹ"���|�����ӱ?_��Εk˓������no�u|�0�HUNzSz�۩�e��V��$����2Z�������G�sxƸ� �%��1��� H�7;���hh�G|��D�#�ת��tj����pÒ�>�E,é`BXF��f�n�[-4#M�6'�)�r�$��u �b 68���Z\��M��M�#�[m�	���?�,��R���'�ySA�8�C��Uu&����z�x�����y�m�7�|�cBϭ])���T���lly�'A[��щ'?���(��+�IT����7ȣ�hm�0�`��.v#Et�k��7��p1�XW����ҙ��s����z��9���MI��g ��� "�M�@X���G��������i�����`L�
Z���E;3W�U�v=g2�(&��@�Y�
6���3w��2�Rq�%��jUW�R�u��R���-�}��(]
�B�(�%G�Z!)(j�ͅv��tƞ1V�X.�^?�D Jr��*�jv����lF���H��z��PF���\W�̼�j�t=�$�Z�"�z��6@p�2l�0�G�w5H�X%��qӟ}V�x5�JP�q�[ő#�zN\)�La^v74�1��>�������As,�}!o���FrϢ38w���+���C���UQ ���>k�~G=RV��Ř
	����5��7k�� \Gb��Txؠ�H�1JR�ڂ�<�a���1hj�&<]���h�A�ՒY�`�8��D��P	`O�9��t�
���Jox,UO�|5�cy�·�{����_�#D�FG�)��z�V���t�V|�c�s�<8��siw�c�po�cc���u���p�1�T�X���{ڼ�gwM���F\[�9<���)��� l�����x0T��H?��6��G� *�f+�7���r.!RQ�� D�z�>�a�z�Ǵj#��Z�1r:)0�)�:�#��d!�q||�
�H!ZЊ1;�1�����-�	����EaU:�u�$��q��F<o�z����X�M���ɱ\{����;r4��_�/w��3E�����b{�v6���'��E�o��I.�i_�k��K��%W/v��j L%�`j�t�z"yLC8��$	�3�Ր��ui]�YE鍂� ��X0�[��t�m9>�į1��L��H��w��¥٥+W�֍$;�QV=yt�>7���ЌǰŤ׹Pd�E�QϥQ�u��?�}��c�VK��$q�k3��I��iǓuA��\�LT� 	�?�Pz��;�]�[=#�$�1�����5�}���?x��	;w�@�D�y2`D��/#�52��ۧ�
����z�aKp��)/��!V�1�VoK�֢f
� �J�d�ǳ!�BX���@���'z,�j[Ҩ�I����h
�Y6�G@2�VjP�5��em��<\�
�~�w��>��Uܨ�P�t���j�
GJ����Td�`�$�@B�� �0�\��ZK?W5��J�Qk1S�v8���h�:� b��uT]��I�����Q�ַ�rR"�yF�Z4��f ď�U"Q:9�aj�����z�s��u�P!	ڣ�ATM�u{�
]������x:�������_ݓ��n �~�KQ���3Do<�ap��~��Α����lqn%9�@)�O����\�d ��(I�Q����y�5�8���b�(Z�o�tA"	�"��!�|�����!����w"�RQP
p�
4o�+��)�"&J}��s2-e�Φ�;ɭt:�#���U+!�g��,)�7��K�8_�a�P�W�#,Y6��T���ږ�,�~}�2��:�6^�;:b7�
8�C��KwsGwԖ��T��e��&�y4���E�qU�_��l<#�,��c5�����0#�e4�g��@���Nj�7����@�q<8օuH�l�7�D�ʛo�.oK��%��Q��"��ᩪњ�h����Ce9�Tfx��F"?]�����UOk��&�NX�,�����A.����x 
��"��C��{�Qs^�p4F���ۧ�X��7`h�;)�S�7Ü��FT��R���3�W��:$��YK�u�N�eqN=��gR���Û)�8�Y  d�F��⨋���V�������T>�{k�%��N2F���~]�6ט^s4�{l��jw�ک1=POs<�KE�K������'j���(��1�5�nU�/���72��i�ɨ �Hh�Ŝ������N��r��Ri�ɳ��?�6B��c��q�)j4;Rk�Hb�3Q��f0Z
ϯ�"��{�^��hDcp�'�e M��k��íI�VF�L�5���*��(y QM�?��
$fS}���R�������z�
���ՠO$De �_JS�5h�6�@K�K(���G�J�/S5ra�����ق2a����p �֜���߾T�u\Mui�x���J�F����K 6��N�&���q�9չ虘\.��[�3��8����,#/IӬ�QT[F��Z#^�>�ʸS�
QHJ�PzM�xT�ʥ�Rg�Q]DSİA��8>��eRm����dN PӬ@MY�� ���W`�Y�3���vAN�5���th) @�ю͍F�po�u�s<R����p$�Ѻ��c�����as�?�����ؾ.�q��B�t&q�.�WnR�x4���s�	"�:���Z�T���^�bl`�����p���\��<S�BpǓ��S��(^=�Z�k��,��/�!N����2��41<{���.o}�X��&�D�&P�]o$F��#�1þ�(���9��j��{'�HB��C[��$�[a{�g!�()�>���b<-RP��<sa�N �N��_��h`���p��E^�������ٱ,��
��@�+��џmdPg�@)KL@���b����Ď�Ӆ��x9�L���*	x�	��0P��7D� R��f���
A�]�j����}��"Vcy��+r��;�<���E^Fr2��5F��2�PF\�+Jue"��'z���* 6)���j�6.���}�(��g��=x�S���H��#[�W�GF�>@�F�����/�Q���l�����WP���c�t�E�V@�I�d]@�(	=�'��A	`H4�-Fc��#��
8bF�P-��_�!M���@A��RdyLЀ�
;�q�}ڣ>�,ӓ����`<@ܢJe��U�>E[5�Ǟ�d8�ql�����U9>9�}��tPlo��R�c��n�Du����*(IzR�G��1���)��÷d4>�N,��v���a��x:�@|���޳�Q��ǃ�؂�7E����
�~\7��O!�D&ė�Ə��A$��u�ID�cs�Y$1�A>�4dȅq\D�@�8ioH����e�+�
�3������	�YT ��>�^�p��R�C�F�,Z(̃g���1�tBF���L�ZLƌZ�:G�v��O�a�X��t��4�al!�����瞓��mܧ��2��m�[����ϵ�����K
@z
�g:�̆:%V:N�G2�$Up\��:�Gz�}�]F�Miɠ6�qt� ����l_�����)Q(O��0E�CѶznj���գ��EEaX$r�RG�mK5z��	TIp)H�}��lm���������ٽ̅��^�F��r��҈`�o�~���<|��Y'�.c ����R�7d� �W�-�
�$w"S��:QN�W�� 4��A�=B�DX�|[a◦e �#PsϺ3�R��C��fs�
%�H9@4	i�٘�&A�D�
:b�&׈)ό���E�[�A
#^�w��(	�ͬc��,Q�j���V�!/��*�h��l����m9>ꓯ�<w2�iX
4�Bޤ���=.z�@\��%�#���tl���w/�J�V���`x�r�z#bI/@A���Ղ2�V��Ez0�v�=�]�����w����[�^���	�%�9��!�d��(G'}6��lut<mI2��T����ॡ׀TYTT��6�|�q�e� w���9�(�j��� f��A�b�{��6��v��}�*+��i�ȏVud\�.j�Pr���鵜(�½������&y���D��P�ֶ䰡��ŗo��vO�ޓ�^P��RW���|������I����k�{
 q�x#:�����RB�
�P*�3�[���6c�,`��D�4�b��(�Fk�S�. c$̒���%��YE`��4r\�ȳ)OS+]-|'��^�aN�~M8�f��^=�|n�F��Ua{ ,�i^�1��[rWTp�
��@Q?T�AxQX̕�����\kv��i���p4�@��<��~�P�|�F� �Zv.���n[���Yx�[_���w����]�u]lJ����WG	�$�!¦������I?H��M/k��E1��p$E~��x���x�����B��N�ª~���ze'.���U������OecW�� �>���ꂍr�H���|S��}�v��$؁0y�RD¨?���.&���'��GI&��.ȧ
&�P��~�L'�d�����It���(�L/�� .)�E���z���kQF\p���X�X'��
��+VNi*�r�m����&�]_c��e���[fDs�i�r.��B{���(�N��\�]��T�=@B�e�yH~�@=�$��I(Ĩ1M&S�{Г�>��M�[�����X�b�:V�;W��BE�߾��k�߉X�wr<�c��yooo�B�`�)�{���[��Uu!?&����q��Upp����i��7L �Ն�mlHth�����翾��* ��ށ���ȟ�#�D@��~g,����'P��,���<�T�e���.y=S�@�)�F�8�i�g>����B��c	���z�Ŀ�~�U+ u Z�A✤􀩧	��Y^�hs����A�n>�0��]_cU���>�)qر>6�D��t�~v�sJ��� ���0�{�t�X�*"S1��ird$
#e�17VC�m�u2�JA�M��e��ATD�	22����v�T3X������Y���X�! �X��К�d@�/��:�}�$��Wt��<!��2-A8����羥l�(�K�x"es�Z�+#���m]�:�-�ڀ�w"���P1}BR6�Hp44����@}]��:nO�B��+��v;��ܶ�g�"�h���1���H�E����_�������n��W�.�L��G��'����{82�.su�"p���u.{^�O�b{j���|6] ���@��_W�F�g����U�쨗��^�o6I�{�`���k��Z8>�8�Ǝ�t����Јh��{G���7����ua����3"�2o�ry�������*I��pԫkSڛf�"4F
af�V`�%/���oх�l�JJ)q�K.(�H�r�Vmb߸��W�oj����҂��EVni�[�T�Ioz2(��y���Aj��XE*!�Y�<x�� @+�b@";��)��j�R��NR�{�?ț������I�3;Q�0�������$�"�\�zI��\���և>�
6��j�H �u��%iF���B����P4�SB]d�77d>�dؿ'���g���ի��+H$%��G����w���׼�`��]���Y�0JS��X=A�z� TeTp0?"pE�=v�kmj$s�Gz�j�@�%ʍzK�NB9T�T �;��rjB�x�4�$S��CG]��;zNc�Y�B�C�����m�01�" "���\��ǼN�α|k��{x�/{{d:�ڭ������5���\�KFR��l�g:�M����Q�>��G=��եZ�%'�"Z��Ԕ���h�[���$��D ��5?ȃ/$�e�Z)�0]�����:�����ƙ۠Ty� yF~
R;3}�+ !DJ�I~S'f�Z/����F'}F�|'��o�%�Fme�8Ϻ�����F�����-�{C쩂h��g
̫��f�c���u �_���ܼuKn�� c J� �V��I︧�"�"1�4������u��~���7_�cp(��T0ܖf5f��˛���
���w�D��q#:��V�����D/��o��X�����<���5��0��>�$�1�4#E�#�u�� �=�|Sn?ߒkW_���c��s����~���ַޤ���چ�����z�/_��x$�,�׫�z���|��?8��ñ~��OM����}�Г__�,;]ݯz�CO����C���F���?S�S�y]]TPږ��k�lf�(~#R�Ee��g}�Ƣ������g�!�DM*Q挈���Rrڑ�Y�'�.���b�"�o�(L�,��I%��لBO���:\��2ͭ�ZfǺ������U Vew[?	�do(�s�My�z��b$�M�(�1}�0���Wd������Ht���w�p_y�e!��]FaN�ޟ���[��:���NkM�WQP�マ䓾���H5���\_��s>��sA
��j��.����SPis��>c������CA"!�bA%9R�b?!�O�l����c����Ciw;����2\�Ě֊_���F$T6[H�t��,9��R��I��5��)Aq��`��|�I+Xi�t��3�> �]���-S�J�g?:!u|p�1�2_�Z�{c��2�UL�61	T���m+ o�|ؓ��	�3Yk*��yr�����p�I�G�Q���$�m+(~UA+jfl�S81/��0���%�Ns���(���Dd��EJ6a��ʄ���cW��Z���uߤ�ťI
�T
�`[Hb���,��� �F�5�3 mF�<�q�*�7����҃�Ñ`�s&��l��^C$RϹm�(�z���1�v��5y��-y�k�����=O�ո~��l��t�o��koT�p�m�U���� �n�~`2^Gӷׯ��t7t�����ui���)��tj-�y����[G�S�5 �W�)����&&W���Dr�=�-� �����~p�ws�r0?��#���5T�W�R:a�����N�C��?��\���ɇ_z�Z�<]@�
 vww�^����o<��߻}��g���I���"��\��?pxx����O|��?{^׀͖�v���w���μ��wX�~���`Kޮ��D�'����uɡX��zC�.��5��>�Sw�N5��S�t�-�4����ΝR�ꆨ�}�����Q�:�y��·N��}'��w���uUe'K�i�����ͷ���u]�P:ԅ�屑#ӑ�2�\�J�z�L�U�w(�?�Z+�g>�U|��,���Tn\���5
pf)s��qS��HM���}�1Fd6�����LK\��#W�n���ܓ�K����Yo��l�,�D%K���)XM�9��	�6ptךL?�0vՖx[����=�W����j��ެ:��l:��~`�4��Y_��k���g����
��:߶��+��B
҃H���+&?�jפ:/�
����|`t�iG������i7�.蚻�k���J ����,x2�F��ė�.�r�H��x�g�Vi0�����pȫI�L��Κ����W|y��ݱ��G�/��T��|�cyw�Dr��	g������#�l��}p���1@��D�_,�W�oq_1���\��}���E -����=����\��K�Q��Mp*`�I�ge�iʿ�Lﰪ<'2C5�>��W3Ҭ��ˊ��+$�z~C&:�rT9�8���1�z���?p���u���hm��;7o���8��u=x������w�z�G�?�c��\}�j|��u�+pg ��s�u�n����
|�T޾7�������&~���,�^D��v�Fy�ɗ�8��6��G���d�O�u:���Tv�k2<�#������}Q��_�y��:�Cy��;$�u۝��}�ӿ����oݺ�_|��1��u]p~���^۹��˯|�o��w����x6����D�zK������?���H�0�4]|�jT$����_�D�џ����Q��t�V�u�4�c��\�H��,�vfj[+k'�]����0	oFl�K���/��8�m��� ��`ȥ�� ����=#ڱaT�ZЋEK$l�qB����hn��M��Fs&�k�\��ʇ?�&��Tc�wBH�:l2-VC���>��2RW�&w���{w=If�G���-5���V���@�ʞ����&����/GÁ�9
�#A�f]:��X=��/���:�ٽ|Y`$�� ��0�]��*a}!�c]�ޑZ=�5�Q�+h�X_��	|`����S���4譸+m�o>+0��=g�\D�@j�H�c�*  ���9ˍ}YS�3�b�73�Pt�ɳݐL�9��:7�8l>���m5f)�|��h2�}��6%���R�I��̈e�{������rN�3�i�P��4���`�FU9�6�Yi��C�&���6�c�s��x3���I!׏a��kx2a��hR���V�w��!������W��~&��m��)�Ա�WU���\���z��Q��I� �I�;Mw3�g�����l*�=i0M|:��(�S��l" q�ܫ��ܾ5��P��P���Q�Nǉڀ��?��WtL�l���>�c/~��\H_^��u��߾~��������>�}��Ik�:V`�M��/|��?�A����t�}o�U!��Q'��۲|_Ϸ��s[�GK��@}�X�'\���{�B�j<�]D��v6���[׹��E�����~ja�E@����ƭvNm�������G��c��77:��������]���/�t���S������_�'����o�[�������|�C��=�Q�xYU������*��t2��W��k	ɓX,*5�-�τ����ڣCN�,v�0��3�/�]T�zi��#m|a�d[,]����S\n}D=K��'B���g����P	�p�}��%��/�5lT�2g����-����ؗ���|�/ȵK#Yo=�N}(�A����yAHUJ`��~U��e�r�1�d'�����H��.��I�sU�6��YR�6ds{KN�D��)Յ�b5ddI�u<ac5���v�4�H�!���yY��g=.����z��.G
2@�k��z����H~=���ٿ$Po�B�'�!���&v:��z�6w��X�	�|U�j��!(��B�WXa"&z�xЏ�kY%�0���@�ז��V11#�zeMz=2
�[IK��� 
����@�8U^/�_=^pL�;D�yw��Ͼ#��Bv����^�G�P!ȕݪ�l�+?�vѸ)�BE�K����L��(����_�$��K�{��+o]�+ jm�ɤ��l�H�5�3E]��(\įX�c,�Cq�3����9=����sg�d��ɺ�����B��`��-1��ؼ*\d�0�vh�o֝AD.U ��5Cg�Pr��4tS����O�{d�@�`�[����_���>�7oܸq"�s��'?�@������~�w0��EX���{�О�r�\���@��L��r����թd
6���ӹ��:I��ܛf�a^lOm�������������@�#��]#��-5l��]�nt����-m����G�}��R�u���ze�o\�z�g_xaw��{���ԗ�ח뷾�����/�{���?�y��k/3�]i4��P�� ���F,��Lfך����Rom�; 	�	$qY#k
�+Ic.�θ�.��<���ԵX���b��"v��Z30�s.���{~�B� %�0��UK��#�2� �r'�+9+)��KT��G�Sj`��o�_�v/��G�����)>�|rW��U�(T�p?Y���$JՐ�b6��Lb^W���T�h�FZ���L�gAV�ْdkW��Q��'�,���K���)��p��X��E�K�5ٮ@�@�z=6� ����E3��(Z�T��zA5T�n%��t4����Ac�I1���H&ɑt��t��*�� �I(��E��
S�k�[2��|П(0��f�h��@#��5�UVB��9��*�	C����	T�|�bh�z���l��+���x�H�F (@pE�0����W6K]��PLK�9'D�o:&^M����2r9��:�<h�֭��"z�#�/)�Tt�֥�u�Nt���n�j\����_߹������7���k_��X�n]_���������5�+����"_M�<�.�r:���)�!�3��g���\j�w�(��n�O�@�}X\�z���%���>�*�*D5Ӊ�(
�R(Gn6"����i�5��m}��/����~��a^� ۧ^z	��g^{�������/}��	���/��߀��Hn=��:N�M�$�e��D�''��e�HNǩ>ι\lOm� �Ȧ��4���K,��.X�\�Q�M�+|Q^�u��a����u[�����/�o?���u���ǿ��~��~���g?����{�~�<țw���C�P:cY�x0�i(왁��d���:q�{#q��&�yfĥ$��k	{v��ڡ再_��w٢չ�~XV[�����9?I�E�$���P�:�:���0r�ç�(�r�@��FE��h�/_���/��������?���y=�Fk��N�{��K�.�"@�A�Pf9�|K��c%���|�I�'R����t[�
r����z^��;�k�]���-o�z���ǖک�s�'"1��P��u��j�5��Q�P,�����v��5�VA�L<�y��W�tI���!�w�1��,���c�Ѩo��U�
�N�m��S'l.8�;0������8 *4LgԪ �Q$S��'��r��@� �dW6�轘��@@��1���j̲^D�Й�WP	1 �@�J�P7����Qѱ\ys<Gc i�ץSI5�)�(�o����4���V��ؽ[xݿ����S/����������Ʒ���������	�z�2MXF�O�2�����z���H�sv�sz��c!��r�����2֕�J�:T���]�X�o2�9���� �(������� �#�o\a�^�����_}���<���k�w��n�?�G�{����#�\ߑ^O��@��nmR@o�=j�3vEI��L�b{j��xF����O���N�h.Wv�re�.z�U�q����0�\�4~�k�ݵk[��|��|�?�'��_����g��`0��ۗv~�����x��o�#F��f�%W�.�|x$=�N���\���lH��2K�����t�!3O�!���e�sO�~��W��i$N�H(����zX��X��ӵ0���X&[dNԫ������}��s�x��mOP���{�#/�G��?��̓��e���$=��~п��b�!�tdM��&�]D�$TＱ�2�	����jm����}�L�'Vj�1�6����ј��˲]���dO����^�]Y[�T�p]z�c�O�>�u(͢��Y�ۖh|�쁂Ȍ��ӆB㶼��!�)�e�8T�Q�uq[���'�I_�s[�J���8^O�Hfi��>s��"	$�d:S��h�Q��TЄ;���E�|��Cq5#��H���
TBW�\GSB��&�+D �:jaS�##D ��D��
��u�E/�	�h���TҠ]y7���P�W7V�G�V'�v������ժRMC��x���2�y0(�R݀��X�P*��-���~w�-j�����zC��������?����/|����8�򚘠�.\7A�9�1c���Q�@~CX%�b�H	4V	�%)t��Y�D��p� m�G���
���$i#&�Gƫ*7���J6%9���,�Fj%R�|mW^|�DU_6�ڿ��G^��n�z]�ۇ�u�^����oμ�����ݔ�`&_��[򡏾,��H��>7m�^/��w'2N	�Y�̍�A�@ϻ���n`���q�R7аL���o�r�ƺ��&W�x�۲��._�ڗ���o��������9�ȟ��Ͽ��ko�y��hԪ?uik���b�MA��M=���>u`�
���*4��u�vy��(��mXU��r�b9�V���ɹ�9/3��-�e֦x.������o�0%1�vW2�}
Ό�obb"�{A�w���n|��/~��~ ?_I�?�fo��$���8��X��p��NҚ� �-�B����NGc�o_���D*՞�R���#V��ǲ����@�_ ��<���?���C��k�w�RoS3e�bO.��ά���zs0������jX����e�ҖC�v�1׬5e�FԻ �ࠪ ���C9:ٗ� �A+Th���I�Eߊ*Ż�v�e��VEҐF��V��X�=A��]@�R�?7o%���(��s��W�8]�?`�����
y7x�V�8fNɶ$D��=ʫS�A��-�]��f6��אj�#GG�$�O�ʕK�~Z�z2�Ҭ�����ZG�uS��1�3�Tye[���_�~�u�/��y��c��?�◾�;�z��'�Z]��jE�ET�E;�W�*��/�"���΂�������p��ѕ�Xp4�F�[V�Y�L�5}F0	�3ӣA$P�1�#:N#�xAs�(X��\cߓv���������v����7�|���6�y���
��<�e�Ֆ�:%�H׵BF��z�W[^��^ ���]��gd�qJY�PG?��tUv6=y��ߕ7�:�f�I"��V�>����;4�-���ge0������x2�1��u�t[X���} ]�Fh��j�Zj4;C/膀<�,^�(y]�4�%wce;U·�^�V�+�d���(�@MR��ˍ�z�[[�܎]��S�k��
R�c]@g��������+�����o'�O�͆����ӯ~���K�Q�)˛������DYUOX�4��n����SX��
k�5�Łn�;w�+;m
#��.t��e�S�^L�kE�.�>6�T�ν�d{���;�z=h�1l�]�`��^O�u�P߯��V��ʓq�?l����P�i�n�z�ۻ����K�wt(��J�P?3�u�>�t>f7��d)�D�Q�}�����2
=�vץ�@eD	|��z�A4W㏾�V�Rĺ�ZC/��@�Se�����UQ'���<wt*�� � �"M�
� �D�PN�cA�cUKw������S�'5>���J��q��=�iq$SoS�ή�ґL�z�L������͏��������I��s}����}�~��!�[�b^a�]�kh[ hc.j�O��e�$�o���,��#~��bx��rz�2p�6�����j��XB�+L��#����`F�c�C5*��;��������V�Q,$��׶����/����+_���v�ƍ�����_��_z^���:�E����/-��I�ֵ����T�?�B½=/[L_lOe{�8�H�ؾ�ձ����n��ZU��7䝷^g����7�N�?�#?�?����.���{��{��ɿ���w~�w?������Q,	����;r������ZT%�E$�f2��
�U�,�+Y�VB�\���pvs9����o�itṭ�%_8'eDE�
� YL�w�����$��j�A�v��@���E�W'���c�?��o\Qإƽ&�ڮ�m�_[�YAi��f�
�����t��*�艢}�!����1�(��	�5��k���Q�����T��BZS4�K�{8�)�	��^�X�Q�$a���lЍ�F�+���* P.��	o "�d�펬�u����d�M�H����5udS�\���!9*hAN�4��סʉ�Ʋ�[Ї�+�3uW�ChNT]��ܺ����j�qPu�Ja_�;_����U@ �UcsS>�:d���9�TndQH�׫-Yo����P�G=F��I�����$B�y}���*������އ��6Z�����������O��} ���'[��znѴ����;�m�eYQ"K��3����,)��a}o��y�|�p�1N�#t�ǳ
ʉe��,�)2�*q�J1�*S�������Z��+�]��q�޼q����_��|����O��g>���k���׏��"��q_��\��H����͊�o�4M�kr�=��	`�h|7�,Iw��©\�rE�Ά�y���cS>��O���L�o\�lW'h�}�C���o����[�Ga��͎z�����^�#(��ӌj��T�S��6��铜�X'�@^F��39�'o��(0>o�u{����b��+sמ;߲�9�:�O�t�.��V+��\�����_)�鿝�G?�y�
�v$�>�ksM=u����a�2�,ծ$~]��z��_��su[�J!�F|I���F}�X[�<����.�<
u����L�4��%�[��:�z�>�6�C���ɓ�@���h�^�DAA)�]Wc^;��LPRK �=�j��(�<�=̄ǝ:"?�r��!��� i�H�gS�%�ꭡ53�}/;c�Bq���� $��[O���w���G�Z�q�}�8�b���>�ZXa��?��W �m4��k�:� ��k䕀���S��Q�Y�f��������ef� �V��ʮ�pgNf�<D7\����~�H	4΀p�w�Z��-�r��BQ�92����zK�,�U�������4;;w��- vw�I�2�=�i2r�J�r��*O�REJR�fUֲ�vي+����R���g�4e<i4�Fӳ�Z���l��������o�9��h�IvH�_7
�[��������8U��v�6K
�j�݋��{H6�hڵ�;A�s����{���_�p��=���3l�`h<��i(��6� H�Z����6�4J�ɩ��31-��ELp%Ï~�Υw-��8���١u���O���/�������Z���]�&�?3	ޕ&��;�C�'Q,\��R�\����!���ܢ n+6�����ȼ�~o��B�͏rI,�L����h�t|/����v�^���(����0F�P�w�y.>@��<�
��9�Puh�֠<��ǟ8���{-*�xD&O�Y0<��F7��e$�ʃ%(��bn�Txi��.�L�9̃���7��58u�X91�&����e��j�<�	���`�/��>�4�%�r���ӦI��8}AD��TCA)**H%ERR�QgC]A4S���(�@Yd��b�R��"�qT�@�6=]�G$�'���d�t\eR����	�ej����`�P=J�S.$�F�Ǯq.�p���ߧ5н��T��6�H�������}+܎D���oEZ��?#&1l�M,R�I*��Se�<��H5�
�i����f�P�ɚ�����<������bv�<sr�s���t�����m���:L(0P��Xtjj �5���4��6H�����/'������e�I�ЄёTo����q8{�,�Y~���?�]��N���2�ٳg_�k���������Z�ّ��J��]���'�ж�
��."Q�0r�{��G:�$�{9H�>�/��~=Ǧ��z��Y2@��f�S.I ,m�%��Sk_��J�I6�J�g��n���]��˚E#֩����n�E���܄���ౣG�o_���<�-���w���1�����t�tk9����z���2�˩V�,����;�TO�d(x�i����\��ĩ
G��<x���O����GD�`�Mڤ�!4���R��(�'L��$�x�I�ƞy��"i!=1Y���5����8�"N`�x��{׉��A��8u�P�,�\I�zJ���	�/D �4E�	o��hˤ����6H"�M)�I���Ҥ���EQ��j�Dk4i��x9;��Q`�*��y�ka+4��Oі$NI� uD�H�^\�))���.�͈7�;���_7 j���P&��4�ԍ��Y�7�}T]���u��f�kS$+p۬��rsF�ڃ�� ��.ᩧ���嵿��p�z�:�z��*��'���:��Zp�s;��@b� �� �z����yR1�avv:�*�C�	��s�����؁˻y��'�/������z}�6@���G�����̀e5ЀS���ʑS�˒g��J��*��q�F�;��	������g��an��<isH	�B�a��IRֺ�7��5DV��}w�=��a�k3T���6d
5[��ʞ*ͅ��D�`��C�an	G����!r�@e����@-�t��9J�B�P'�
חn�Y��	����I_�)��'��9�H������t�tZ��Y�m��ыN��k�9�  GYh0���E��A����E9�v"(DX�@�'��y�D
�4�Դ�AlmOȊ�qO/��	��pڅ�����m�}�y��;��cW��^c�r���ld��/f�(���F���*~f��!�8�Rqp�v�J68eJȺ�yw��4V%1��W�r<�5#j�������n�
m�5��Z/����IJ6�9+�E�M���p�t�ID]T���%Nk92M���w�B�ѱ<�,�ѣ�W:��"fg'�狅?,:����#���q�������Ļ #�I6�
p&#��T��W���ظ	���ѱ���6vu���X�7���.V*�O	/,���e8z�4hCqC�aW�����2n���X4�-��q��ś�:^ݸ642�C5U�\dq}e�}σ��S��8J2��Y�>u��[\�@�9T7���Ba�5�9�#5X�xԭ�9�!O&n&-�9�y&��J�Öo6��t�q`rb?�Wp�'I{sTa��2"X�ǭU�02��ri�C��NI���q�r+�k4��Gt;��#ǍՋ�;9�?B��N�Sa�w��Z��L�8N<]�O��Pd�y�D\�|'�5R�/�FBA��3;��j��q"�e9qH�	JJ��A�c'�A�m|���m�		]OlԴ=��)jAC3O^̧�q����u<>>�S-�sD�b���64[5(&@��	��0L�Uo=�]C��Ąj>4op�Z{�k;�0��v7�F�����3�
�H�����N�p�z��S����e����8�H�S���RQ��O�WO��~Le�AF�(�~1W�R)D2HLndpN�>'����}�F�8Na'1::�����K/����l�j�:�#p���е�֕����dc� Q�	�Q�ce��� ���B����T��r�]�kw
'O���������5܀�b�z�C�n+<GBKg:�}T�m*MVoC_���u�| dέЯҘ�;��ȼ=*��&�RQ#u8�qn�;xog���m^�g����D��::z�2��s��1�n4ڠ���N��`�	.�����.Lэ���&�0�o
L��vVo܄j������B�ð�����3�t�"�U�ٺ.��(�9�062�}޹�yܢ�䳉dd��# �ب��C'UR��ꀇ�����fR�m��1���K�6�=H�8�Ld���v�K~  9�IDAT��|�>9n!�$G�����B<�����N���hJj�t�&yl��Y�R����:)u�㹠w�c���y-f���HC��h��	��R�q���vI�A�.��� q�A�;,ͯ�Ԏ�9�*ZD��hܽj:���H�u�Z�<���ꬽ�͈��[o�>٪zk]��h7Aƕt2sJ���&��ϳ4hҋl$��NŽ���EB��"��A7I
��B!�����T�ַ�O�:�V�\�אm*<�&X����m�${�m����'GEu��(�!�(�"��������"%��a��LC�D.�ZA�]68�IQ!]X�	h$�r��cbs�^Mx�����-j2��n��j�jg2ʩ@�Q�d��֋�/�U��I�H�y� HIJ:*Sm �]t� r��7׼��
���n�7ށ7���� �I������p��R`tf?�+k��K]$>�`n�F2p	�]z�ŸF�����q.�\�F�
�#eȢ8���i��W��]��wJ98�^��k�|��
x�����<�nZ�I�%1���#�v!0l�r�G��p4$g�SAQ���E�)~��V��G�.�uEj8B�g'!��u��ĄOc$�²9�ĺ4!ǯ�"Ҙ���t�� �B�#��N�IS���4r��7p��E�O�>>�&����	`����5,��Q,��4�O����]���b��Q�V�T��ڈ���ق�
�UD�zj�}���i}���"�?⍿�/���E䃩E,ļ��U�ۖC������D���.}.��
������ӻ�49v���1�~c�בUP��-���[:�� Hl$��#��ׇ跪�\t�E�A�K�����̉eo����mu5*V�����e@]
@�<���ȱ@mD�T�IG��+km���-xYd��"[q���i���)[<A��lK����)O��4��c�<��t�f�մ6z�fD���g��w�C�;+r�U�\�	k7W��|��4�>ǲ�.	e:#1h5k��z`\Li�U�T �I��ʩ�@����|ܘ���\�$FBbT���m�Xz�<s�d	C
k�H�"i:�w��w7�����
kp���FY����0�,d�$�_�v"T��bf}�"��3��6��P�@)�|.'�����H<�ײ���u�$)�U�CD�����$M	�F
���ګ��p�	�<�H$UM�D����Ph�u�֠8X�.��#�Ƀ�d��R�|�^�U�T9�4>6Tl�w]n�������)�qPBIӒ��_ڏ��G`c&I6mVI��ޫ�J�YN%N5SD
�#Q��<tP���u�< 
����n.//�E��sGd�x�%�ںB3�Hׅ���H<m� :ݖ��FH��G��F#��Q�m���̎C.g�BG�.�]]�CCC�R� �R󥼸��(f��7>*����E��YT�W>A��Lk#C_m���ԭ��ߊp��3z���,J�Wj���F��<���b�<m�W��~Oup�A�`��\ŉ��=\ɅFS\��ɓh��<��G#7w}�n�������3��?��c<��lhyԊY��Z����"n�jD�Y��q/]A�1����Q{"��(L����K�y�y�Z��8����NTW��(����*o洱s*�6r5-R$�j�JP+i6&��t������qj��ج4-�}�W/F����uxS&��Zb�����͠�j��9��X�B�fῃ��|qu��\�@��(��so��uA3S�}[Hʐ�p��S�B�Bq�P=2&�VT�e�k�M=7����_y�Zh�q��= ��OƤ����<e���e��H������wJ�d����ȕ�y*���i�ݿg�%��+�4e�N��0��R�הmkPk4��[��&`��Eѝo���0l��<��5tp9�
IꋙN��s�0A��=UA�	�[��r�g�|ܤ�b��Qk�\w��z��<N��'KCe�L���*��1��Ƽ)w�7V��4�����2�1�f�7�#��(H�(��\sq� ��<�[akT#'��&�ipo� 5�ՠ�.z>�n��m��`�}Ѭ8��kOᆾ�铦��D/��o��k�+-��*`t�(��Ꜫ�7�x�� _@�#�!"<j��.ڤ�xU5*vd݋���C�����+19�yF	pB�02�.�?Hř��9܀�8���j�\$jo:ul���8�.FhhZ�F��vy�SU����k#oSbò"U)R���2�ix���#Y�G ����c�(��㜙�P��!��!��F
���j�E�[x	K[j��p*���S*�aǸ!Ft���'�K��X�*	jP��ۊ���5d7�Y�=ǯ�ͷ�8�Ritp^תI\�BEh����N��N�T���)J~1Co-�72��������A\�ꦵ��9YƑ��$�ɢ�\@��+��cbX(p7�ؠ	�&ѹRNQ(���$��\�djE��#�4�H��)��F�Kl�${�m7�zOL��}X][����B�٤�����Q���n#!�K_��'fffa�Nt��̛�y:HB"��
�nQD:4�<����41��(�W߫� ��X!����H4�"Y�Z�;��ò�I����vcs�����z�< K̠Ȇaq�=}%�Dѣ��BJ7(l'vwV�΂?C�?w%I~���̟���e�blG�᮫J2���;��2J���W�a2�������O�a�`������oy<��u��V�� �`�д�>���Rue�$,i��Hm��<��9N��+����Gq��w�v�0��� �rg��Π��g�#I,E3k�atc%�!�l���s��FCg%
����MLS���i7O����8��T�(�0m=�]=g �P�.��.^BI�/�\b*��(���ja��,�������l�$�E���B��ql���#�P#$X�x-B���;�㹈*�ISm���iV��{n[�L�)��!�i�jO	&۰!�P��Db�0��6�G��<o)��/�%dD"�}J�W�a�}6���D�����1���^*��:��L�R'����a}mIk33����g�^��	|���.��իC����9�5Aj>w+�<=�jB�N�S|DJ�Qŝ���l���
�����cFG'�0�^_��h��,��T�C/��ko׈�+W�L]x��Gk��H0F�'��cG��R~3@"��L��nڸI�<�����Vq���ӷ�۸çxo��}��=N;��]�{o5�RYa����Ȱ��;�n9w��(ʯ�K.�?�D�6_*O]}.�k�U"$U�.Bj,O39���Rv΄��q+4ڶ�s&��R�B34�f�F7Զe�-��۪�����0�M[��4c5g媅B���_?c���$q��!3�</ğ_�?r�}�X��0?�|�C)mDH�R��^�4�x+�ۮ��k��h?����}7^��9P�֘��
�&']�zj�N�4�A��oՅ�rZJ��v���\�p���;8�� P����	J�L�"n��Y0\jö�f��=���{^�wf'�l��7ՠڇ��W��؉�!��x���>�4�g���xY��t��]ùs��̵�œq����<8Kp���Щ���v�����4�W�N9���Jӌ�X�1�2��'�Z�C���-C|[;�n��u��IO� ��ޙAm�j����@}KQ�m�z��f���o����W�p��՞�j�k]�N�Gd	��Z` �(��QB?%0�7+����t�eYf��+�:�z1?���P��i�7Ѹ�ps�!����G�J���S����u�IZ��m��#�	����\�t+b���\��شtb!��k!#��"���ިW��wfR(:�R��ՠ��xb�/���x��ס�Z����0�g���>9^����-��{�eہ����j�>5>>��z�³[ȁ
�&4��~���g)��H��G`����xP��Г��ُ=��E�Ѓ��j4�n6�~<{��onnu����7�R:���+��[o���Ehv:^���D���Ba�M�B'T'��AO���^�*m�1OcUX�߃J�2�-����� Q���� 4CO��z)����C�N���/�#[���1�N�&Ѷ���/�|�R���ڿ��֏j�[�=O/�E�C�(�C�������O�����Zv���k��wCU�K��U�J7��3�<�����E��&\C/\<���&iki�z� Qګ��4/�o�J���@���J起��Ěcҡ��O��oz�����Φ+R��nJ����-C�\T�`���Bj,
W��`ie�睢�=|��:���������?�0??7�ةP+��+P�P OY�jӇEj�D��m�CI6v ݴ�1P��A�o���@y|����2\~�m�_p�'@o�<n��ԩS��<�����VnT�&���*��W��[021�_|h�P�C�����u���j��x�����ɱB���E���VS�.�C�c�7ɣ��C�~�jmF!��	�\��,z�>�'f$:��P�D%��BH{��SJU� *umt�`*]?�m�T�,[k�v�gΜ1�Q������ ��;!�ۚn�	�CQ�����;Kh�d�\E$/��AjE��*<i5UfMOPV^ݛ���ΔH{H��;��T!�Y�k܋pd�R�Ͷ/z�Ws�E�@�Rxt;�o���U��֛03U��o�����p	</�fmuz���_.--�<55��	�^��3��Lix�O�B�6��/���!��������:x4��.����Ì��l<�Jsl#_����o��O|t��ʉq��Nβ�R�E���+�N�|�ݷ�}H���ھ�����z��*�v�O}��"YX^ႲX��XNQ�R*	�*��u�5bQ�ƽ��$�8ӻP2#��L���Z�D��	#�l���鬓(�GG�=;1��k,�EYc �tZ";I:���H��"��,����[ʨ<tD��Zq�^�y��'�1�]c�>�es��#�qT�����F52���%����H�l}�h�~�ke5M��8t"��Ģ���d�t͂�E�8����^�+k���g�]�������Qt��U�K��{�ō�7fN?�i�+++��{��i�\_k@�M$m���v�I�J�� b��'uHͰ��K������CH6����?�!�$pm�
\��z���3}~���g�ø��ߞ;x�����;/����$�MN����s{�ǡZ������$�"MaY&���1�h�)�lo(��T�Y�� B�l\�lb6;eK �G��!��k9��l$���0�Yx�W�����zt�\lz\��tH$����t�.����R�CA��6^8m�������n̊�MGL�I�E��TxN�TE)�@3z"E�n'W���}���xs�cc�l�*���1|\��t<.��
��y��7�jP*�`�\YǍ�+ܝR��<����o�#�Yw-��Aq�s?�ƹW�Rq���a����p��'��8ͯ5��eX�t���(B���F�N&��A�LF��s45�K��04���Fp���\Z�
σs.��Cӗ����{jJ�1	���_;�����?ZX\��$m=15����013	O|�	���G�� U�q�.[U��T�H�H%���D�HrZ��jEd!J�v��0�d��� �K��H��FXXM6"J�>��Q6=�����Bb��"�E"T%��b�FI=����#���w|�B�U�au�����
H�03☇�� �Ll��������� I��J�w��w��~k٪�+ �$�倪��6�Y���v]���"�R֡Z[�f���A������T�������Z������+�����������Z>x��w
�+:��G���`���0�P�3p��#}��C<L�dc�ZS���}O�hN�f��V`f�8�	��e(�64�6�C��*��W��߅��v+�E��~�w��s�k��{�qce�G����`i ����ީ����g����� �p�&��L�u��7-�6�l`A�Zp][�D��"D	ln	�T/^%�����b�#���p*�s���i�9}�m� ����U�F\D����|�U�^����ȩ5.P�!��ƴZ\��z�Z�w*���ϵET�A�D��3�6����c�q��Q�9�H�b#�!"�YM���@��A��k
+���z�_LkV�� ������������4�-�*uH�-><5���T�o�˓o�6�ҥc�����������*i�<�Gx���cp���9{�[1�vH%.[�m�${�=�z-m�V]n�X���a8�?�A)o�P1�1x���չ��}��ĝ�����533Sݮ�y�ŗ?�;_�ү_x��O�(ᢴ��R]���%�؏
~���i��_�
\�r��>K�@�$]���v����X�R-`}H���������rʷ����Yd� z��n��'�#�o��Ű5J�d7GJ�Zv!˭�zTkBF��EM"�{�nZ���]$�՛�J)H����c�^V�L�T�F��aE
y���i�ݪ	�/JJ*���'b���j����/2�xT�Md�'��1�W��Vj0݆}�tJBpl:^ K`;X�y��O���?�y}���;�l�x����~�;����E�W������ɓ016�	�>
�.���Yx��Mpr�"$~�h�Ķ�#c���"X$��9Dn�F5x��

�a�� ��=�*(HJ�E�p��X����ƚ7�x��O-h	���ҿ����W���o����'���G�"aР<2
��-��O¿�s��;���Y�v�'?��=b��	$�C�܈�BS4�3�L�S4�*<E�u���禷��G���W���2��f�1�^�gh{�����fZJ�Ȥ�UnS��m�����	�{���a�r�I�%��hM*<�QW��$\�)�]���S;iD���s<�n+z��6�hse��f�`~r��x.J��R�"���uA�d���Q�A$	��vl���,�W..Be������ځ��z��/��W&&>�f��[�~��������_m��`ك0�� L�O���app���7߅���A�Mɟ�Pbh�2z����dc{h��F4�it�i6�#\����Z���]�O~�8Fm��F��ĩS�8� KsסRm���?��j���{����������k7��,-~�W_�[Q�=~�4��>�O�F��7o���>x����q-��7^��E*n+�Wk �Vb5DPY>;Hǅgõ�B��M����PHMzz�u�E=�VS17��~�0H�Sg3��L� �;r�I����JC���Q�AF��2q�8�m �8�.���H�=�#7�5�f��B�'�r�(k�P�֊ʪ1|?]��ɕ�k��~ְ�ɖ������5�ω{���B�����K�q�!�k%��hV��z�69S^�%�Ɗ0=sƆ-���.,/�B�vn,�=~�ҵ/~�Ǟ��7n�㉉���z��_�2{��s����_�ҕ+�OдdHt(��8PB�چ��A��~�����u�����=|TEF/���`>�4a{@�S�H��:4������A�����uȯ���� S���8��	��ch���*�}��sW.>~p��7��k��'O�Z.�[��ZC�q�6�J�2�87��o����k��ڏ�GO��5?���յ*���S��U�*L�L�������o�˯^��Db=q�^��U�#��	y�7��R]%�����CI<(�ް)2�Q�A��t\uj�@N� ��b���	yd��RAF/���~Ju�\
AGQ(H#��2��"b�N����lt+��H&H��)\W��K�;,���U�!���#!��n7E��&�i)1�k���(�(-�Z(Z[�"���'��.�$%Й~G�%���Y
�ѵ1�6�|�1q_Dp�=h��;D�Cq;�_�G�6A��¤�C���z
����k��=c�P]����
�C�V�!������+G^9��7���/9v��\��0==P��y]XXpZ�����������hqi�i��8���
< �O�4O�X0}�q��؂���ᕷ�������8�	��j}����T�`��~��BhhD.\�9��
��/����ai��W��Sǎ�ؾqНh����۪���曟>��K?y����vjutd��w���w̜�\,Wۮ[�p��OTV�'?�O�x���j�ڄ�l>�X	��u(5a��~X�ބ���pea�x�Ǡ�����~~��y���N|�ś;U�g��0t�Fq{U"��QO�F���Aˌ"�d*���H���A����
��d2��&�d"�R!��	�,a�0�H����w!����w
����nФ[�Y�n�F�mѬ���W��B�'��"�&Xjw��)��T%k妺��I:�d"[���h����V���H�;�M])�	�@Mg���5�6JK�l�5��sI�P���i�x�ͯ��6b�)���ҩ:՞�H�Th�H���V .]]�F;�������å+���?z�񉉱�st|lyzf����?����ɗ�Y0���6h�K+�������gοu���,���)>�����xF��8X�}����,�uU���?��;�T�so���!B;���]�.�t,�f�${U�a.Vi��ţ�}����hvC��3��}����B�ۀ�K+��>�i��A��P����um����W��[���SO=��ŚeY텹y�^,S����<�>����h���u�����K��PEO�k�������������z"�ą\��ސU��(	G,�8�96_i�P/c�9�zQ�&���H��D$5�S(c6�I���Z�3�
����6�5C����/D�8��N�'QOL,Lm�hz����UE���D�8�z�4M�ݯ��Ĵ#\�!���Z��{D�=�+��B*���yAWLUU7�����I4���M��k&���!JJR�Aͺ_���Js�:�$ޠ�Ykx_�8��_���ʎ�D�T������ u���Hb���k��
�ZC+�6�R0�CC��#=˰`hxZ�.,^_ABrm����&�����3��rH�"4_Gu
�f��{	8�����33�v�pce�x;�10<�9�fO�����^���\� � ~/yPL��f@� ��d�\z�Z_w3� ��@�]�\�آ�҆�ߎ�`�js^~sN�����@u:��(�As,�O7p���'!������Ծ���X��tK�g��S���ӏ?���@i�C������"\����g>�<�"���5x��`���B/�s4��-1H
-�6PQ��dC/@I�ZIÂ	�ĉ��(-���lB#�Q��l��JO0@Q7��8p�CK��X��B��9q��u���M�VKGxǩ�M��L��4���(�#�4���k�r$$��c��������f�e㵅�l����qp�8_�q$�)iW��l�D(��T�
ک}$]3R���	"ajZK�A%�.�e�K䵔QQ��#/$r�B||��(�x�j$E^EU��GGI�� a��D=p�6�6"14�YQre&+&:/!3021F����-�����Q�،�V���Z�|�q��wt�5�� ��e$h�V7*+�����`l�,���?|���g`�Fb#�q���ɕI:@��nɚ�m�${ ��99��r��Ȱ���b-P�w�`���v����p��(<qr
F!ɨ�C�QԹw]CϾ���ڀ�ZL�S�!�w`f�x��g!�|��\^���U��$�x��z�b�s0:}�8�?|�<��$k�8.zaՑ[:�;QS�B��'C���8�9�(VR�
j��!�DC��#H�Sx�S�se�b�w\c�Q$Jޓa
�Ie�1�ʦh���I�`da�,]CDF��DhD TM�`� ���MA1�ԛ��K��̦4D�Mu<�)���Eg"v��<wq]5�z�P�l��[J�-=���]\k*Ӌ����t6������c9j�i����Hto1��H��K�@o-g5�{�bc�6��}�ҏ�hqO� ������k��:#�\���x:K��LM� @Gۑ�Utbjx8!ڴ���z�M'''a��!h4�1�T[����ڲȏ�B'���咒�`f�����Y�s����_�����Յ�Fi�v��=$8X9B�a7F;��|i;�c�(B��=�� ���Cݠ�%�	UV��k1y�5U��T�>�yq��D��q�-��I������S������`#qX����þ�	(Aix�kp�9(X�7�'���^(Ä5��M��߀o>O���F����H�pA�Q�-�;���ӄ
��TM"�Y��@nҬt�dZZ�A� -������HH��zH�A�����޴(f2C`C�_MҢ7`Ù��x�dz�a���p�!
��?�E����x�9�1�������c�6���N͗kG�a8F��zD�J�(q��Zй��,���F=H%�)���M���{���b�"�wv9f��w�����,��LS��>Q�WC��%�KѤ`�B�BE2EQ�pZ� �S���/TҞ0�rX�
����� ���SS��`ф���L
Y� �緡��W���O��C��atd���:.4[G&'�¡c�C��+o/�Ko^��O�����5���L����D�<�,�@b�\I4��`�$�n'q�Jx��q#O"��M����5��\n ���{w������e8zd�E$JE�
95 ���|j�
4�UX�9G���qZ-l��J�B�bl�-����v.]�ÍUb��`��lt|���\/�a��c�9:��1HP��+j�(����D��*�r��$I�)� �D䄢VNR�~#�aL��DdAQ{FR�B����F�&eRv;��h
ՙP��в�µ!���
ژ�ة�Ɵ�r,P�iT �ʚ�{F�Fa�$ARD�s�aN����zR�Td�F��pD!�zd#
�T�W�6r&�z�5�2-�'�[,��?w����S�S���=�5����45��4��j��\O�G2�v͠�����<P�T�H"�V��#|'t�s��Ի.mƦ�abr��2��W���X�݄���P��B�GS�i�Z^7�ot�b�,�,þ����S� Q����>�9{���+P�{��6 ���7)
�K"�;�|"�>
D6(�ƞ��!���1�n� �� ]0���..�1�iR�@�Vs�x>n��
���i�{ih��K���9XY���P�G9�?&?#����H��G9���k�HDB��}h�����޽z�<7�$�W�00<S3��ƠV���P��<�.����ES�(I��P&嚩��H��q��t��dP�YZ�l����ygF�Z_y8�j95T�o����eR\����>r�ŕ�����9��6�}g�4l����ِS�
�*��4�����%`�D�Z�miK�{�I�Mh��6���jl��Q�4��!�7p-��RYr��R�HQ?��\��(C�~�t�ODg��P��&��)H�#E�v ׬�ץob{"��q�#��Jr�1@�g�B	3�0!�o-��*�c?��К�K���k�$�&��L�w�ǵ]�NΞ�k�98rh����}hӎ�#'O��1:7����zP*����T'����f��Mx���v^y}�j>J'pڈ":��x^ɩ	9j���H$<C��z��=-�� �${�����]\\�2��yS�@}����%����
4]466n�WV�������F���`&F�<�K�!��p�������y|�
�H4;�TC��ކ�U�7:��h�ä�J��
�ObU�vk���l�/���� D�m����!�qS�<��p�(j�HD��R [�d\�B�^�q��P�X����� �D����������"4�-��I�`��$5⚈nP��r@)�q���Ca�������^^����쳧N�Ȇ�=�����������E���$^ܵ����׮�(E)T*��(i���K���7\��i���$�&(J�y��n3���("�k_G���c�#!��EbM��t�4�B"}h'X�/�5Fą~D�rc}1�R�"(a�i���m��[U_���5Wp p;b��C��@[�å+|��`vf�����~�=��$�Q��|s�v���ʃ]|���*�{y�����T�F1�d؅DI��8�<�������?��0a���V�&PC���:�[��I6�N��~����oTj�l���c�ݵF�f�U���cJp�wL=��걬v�>�%]MbCU�XM�$���n��_s�˖	z�6
I%��<Y��z}���햫�~�Wt���Ɂ�����iZ���$��H�������Iԉ�С҆�Hp)�I���a:]�`��7�T\ϵM�L+���A�Qy�i�I�X�����P(WKhfl��A�Ufl,)6L9�N��oR!g�u�Q��fh����;1�$Ad%���������@�����B��܂�v�3��E,��0�P$*���aǍl��J�j��A�ٖ�p��������mꑅ��0�����'���M���@���������'�a��^V�HXݮ�4;��"��4�=x=�b=�O
à�q@Y��r�a�P�z$���h�A(t���$%14��&@�z�P����e�O���(���B.����:1B��;��p_�����1	�r���'�cZۇ(�p�HF<\(�Xh0�(MUG�`PM�ZҤ`&<zH�5�E�r�����5��M]7,[���Fൕ՛��j��9�
]u��uC�S�a���Z�u�HsǊeuzbfHќ�'�skU��Z���#�PMmX�5�W�j�����l��kZ��y�T�o䔉3�?�կ��va3�x�< ����$����$�N����}2x	�#G �.���+�<�4����c���������� ���+���8��:���I�����f�sL��f3�u�fX.n�jQi���&����v#��8���ۊ�F���8�ٞ�f}q�t��4��d�h��pzq�����w�G�*�o���k%�%7�h��]ˀZt��Nн6��`�.zQL�]۠�vlw|-*�J����������?7OO�یkJE[�9Ϊյuf2���w.7�ݙ���h��(��ɯ�7GG]Z��E��ΜI�g�Q���_%��(�mF��5b�`�Ӂ8,�1ЅhYe�!�r9P+��$�ݪQ���G��O#�Z^^v���B�Ж��t�΃j�����4�z�H\.�i�N'�uR����;*�UԜ��p�������8�pT�c��FNk)J�xV@v�,�ȎJ[���L6��������Z��1�>�'O� �ߙH�NL3��'�e`����w�G�ߝr�K<�؁�?%	��~k��t�7�4������l͝R�[�n'��/��3�J�ʹ�	2�"!��kA@}���x !Ɇ�������hHHH<��dCBBBBBBbG!Ɇ������ĎbO����������)��]vO�I4$$$$$$v
��ݓdCBBBB�a��W?�dCBBBBb�!�ƣI6$$$$$$$v�lHHHHH<��c�$ِ����x$!����$��S�.!Ɇ������$w	I6$$$$$$$v�lHHHHHHHl;��l�lHHH<�ص�Y� ���
�dCBB��Ů���hH<Z�dCBBBBBBbG!Ɇ�����L�HH�-$ِ����@�DCB�n!Ɇ�ć��p%> �#�@��i($;w�K�!��r%H��a ��C^b�ِ��v�KHHH<Lxpb�{�l�Mp�!ϱ����ÄǤ��!!!!!������%v�lHHHHH�8$�x�!Ɇ������ĎB�						��$��������}H[|? �ƮA^��i��$ِ�������QH�!!!!!!!���dCBBBBBBbGqOdc[�hdM�-!%�-��[BB�Q�=��m��Ҽ�r�y� �o		�G2�"!!!!!!���dC⑄L_HHHH�?H�!�HB			��I6$$� d�EBB�a�${�h�=$1��m���;�dC�<	�� ��B�DCb�!/�;�dC�<�G;�A��-�����L�HHl�l������x�q�Ȇ̃JHHHHHHln_�!���m�HHHH�A:�2�"� כ���
�J��h|8<�dC.���]HH<��kXb'����0��"�߅����ĭ����|� C�;I6"HB�s$$$!<&o�ƃpz$H��ꁂ���px�.����HHH�4$ѐ�x�!�(d�HBBBBboA����hHHHHH�-H�!�PB�HHHH�H�!�PB			��I6$$$$v��J�ц$;I4$m��f�U�岀�    IEND�B`�PK
      RZ�7.-c&  c&  /   images/0291db46-fb1c-4fc7-8f6c-e1e807286f19.png�PNG

   IHDR   d   U   ��A\   	pHYs  �  ��+  &IDATx��}	�]U��w����jOR�S��l�E�긴�6��lm�m��8Ӷ��i�eF�3���.�������
�
��H�JUR۫�����sνｪJ�R/����{��{�o��Yb�����;c�SNW=�-�����趍%1�D��&��2�~T�bH���COVf&c\��S��wj!��,�����gZp�Đ'��>�Meҗ�
\W�D!ęжǢ,ļEr���T���B��e=�ʙ�����9�~=����X����d��'C{b��E���~�w����w��W���lW@(p�@-b�u��l�a�1���X2B�%`�o@C�I��Q����o �I��1�u���,f����c`�LH-����I��o���p����� ľxY2>���I<ׁH��>p��uBl?��C������<|wK�}�=w��)�mc�H����h]���8\8���0d�r�Ï�{����n�B�
�����;a��]pV� |wW�^��� �|���ֶZ��%|5��@�5��H|� � �#2x=�սf�T�,��H/���w"|�+Ƃ��������&��=�
}O����n۳�o����M|w����x�e���a�`�|�[8Ƣ%�sr��d,��7�D���H���{ۅ/{��+�]{Y#.�·��Yv����(�ï�X(�\4c�#����E(PCʸ�"�c}d�"�3!��bs��R�Q�f�F�\�EA�K2�Wl�$��7�f /J`�%ij�2�b�%V�G�@�ש
�_���d��o�K�XN��z+Ƨl?�¨7B�`�2t���X��Y}k�d�5Y)��<�(����?R��Wx/�w�������zg��u�os��ղ�k����@Z�����2���#-��C*!��a��[�{ԄH�h�$�g�B�&�&�AS�9�񀡔��1�I���Gi�<���$i6�_2�T�7�]��#e"e$��<j^���PBs)a������Yp�=�3���]�Ҧ����tӰ��5C�J��Q�W
��G������_ſ*U�<TκV<va���y�֦ݕ2*
v	�AK��29(�(��N6�D��#��J�a��6=���}�`7kp��������G&:h%�y�U�B�� m>J�kA�q�ú3�A�rU����V0d�v%
�F=�$ G����8p���OW�W9��Fy+����cQ*z���ٽ�z����a���Ga3
Dn�m^��+��ج�����KuT�7�|K=<��ѱ�9�ɢ �%X}B�G�����.1�Ҋ?�Ö1:w��zزa�������xɥ[��˟�����a��a�!����M7�
����ȁM#����}>|�o����0e6��e2愘B"B2�]�AF�"�5�
l��Շ��o_��O|!�C�t���o�x�p0��?)�8n��O֮��4�nʑ�7�󓙩C8k�zt~� ����]x׻�z���q��n���+��le�$j�Hr�Z�h���X����X~��_��%��Č��Z}>��o@��J�������އ��#1�x���cpxt]�<�� ��4Q�^� �O����i���(iNÆ֬,�߿��b�+��]
=n^�����+7�5t��P��ltÐn�Y�?�(���|{*7;U��ơ�����?�z�9���{1�˕!>������B;d�	1eL��T3�A�.Hj��r!ͺw��nmz�� ds2�8>�D ���*���ݰz]?��~4�>�g���!SB�|�5@06�!�%��'�� 
�㖡���{�_�3�-2�tγ�Y�}w�&�	�wÐn��P�@��.d3G'��<65v���05�f�Ⱥ��#�����
8�H9\r����ɘk�E#,�Y�%��*2e*��"��4� >g�W!<-@e�0�{���B��(��O��q�m�>@��M�ݏ.�����.aӖ��Nq�FC"HdT�E `z:�������S?=��	���7�����W�989���L&ڳw\��Ǐ!�=��
~������0��s3��X�Qb�+��\��ga���:�� 9J���ըu�D�QF�K)��z�;-�!���{?<��a�X��4]P���l��|��؄����n^�%��;G�L����
��qQf ���SVU�xD���6e����G���}��+~��Jam"k�?��oU�~�G_@�����ǐZ����;��=c8Hg�h}������o��98v����G�1�L�$4�0V(��1����W��`p��vÊ>X��{��!k���C��mt�ܭ�a�c0�>���8�`��~������`V���­k�Бc�˞�ܱn��N�9س�,ӧ��2D0�_��}$�e���G|�������x�٫/_1�b�[bŁ��������Ⱥ��h���� ��=���N�!��쀜�88����i$f�f��߬Yd�������8���0f������T�W�%��i�D�c�>^��i~q���5�Y�q����"�FkU��� ��={w+�Tp���0:z:x���t#LO��԰�::��I4ey�FԱ�����t�e�P��p�-����f�������cSM�q��޳���L���0}���������4/@-��50��OB���É�M�1x�KK�\1�T�}�g �AmRB.Z�4#pe�� @� �AI|4B&�P�J&�)��ӽ���S���#�-:�;�z-p-�B=b��50� 3�����?ډw��ɮmA1G1��%ş�Qm :▥4�zl3�]�Ĩm�� ��dПEP#��������kad�z�ų����!�޺�D�ˈ����q�8�\���l����-C��6�a���#�'`��J�h$s��I��aˈ���|3��L���u�Jg����c�94>i.�?_�r�4N2f�,S�QP��2CXg�̣ԁh�uY&[ �D��d��^�03��i�Hn�P��A�X��_����{]L�`�3M#�����]�A�5e.��!�
�@ǅ ���q�J�R/�`5a����d LGW�2@�K�=2�pE0�"7�{�.��2H1E?#sunn����:�ef.1�"��}���i�'�I�N��kW�<�Ь����Q�m�"�M9��jǁ��z��R-� H2�t͐�H��1��cdz�$�ԺLrE��`����h*#&��"��Km���0H1�b�T���.���A�E���n_3Z�]]7�BƦK�/Z��w�v��1Bp/U��Z�2GuU�RQƕpiTI}A\*O�t�"���$���#��3��Fc����:o#ng"�m����d��]�����i�q�%&L�T��e�ni���A	��_HCX�������?1� :��z��堉̢G`��Dg�|"G�ȥ+��>�)]3$
�LXJ��H��&X�� �y��X���g�.�4rڱr�h�LR ���8-����X�6��U��D���EdZ�:����qr��P�m7!���$�.�/ʙ�t*��-�HLܓL����b�\�vD\���>AYXJZ�JrL��v~N��	����!h_�5�C�Tι6C:e"۪���J� M?i�*��H`bL��G��!��g�NVP��0��uB��cȩ浲Y��l@6_�ͺ�8�/�%I��DMޅ�ХL�m&F����1�&�c`��D3�t��mkA]�� b����� EJ�G0ĦTO��ƷK���S�3*�����c���J�&+�U�8��e3c�ʋ���D5ӊ w��F�-�ӺU�L��"S�m�x��)���m�j�obָ�&Z&�􋩄$�|���B<�f�eЇ�d��"r��4g�x=��!iO�R���2,3�F�lb�s�>S��I��?���n�Q�ͳ��FZ[ը��AJ�.C�V��)�O���qi�-��<��eP������`��S��4��d�,z;Y��q���oQ�Ohy�֐f���<ԛ#�<�~��	��F�v?qȠN�`��1���@������l����n�lڦ�Љ��YO�J�o3�T(fP�M#B���L�M�{P~�����;^�io��u]v�US�a.,NH�y9ռV�rU0�"�b�-�8�E�m�X;Iɷ~K��'�������?2�.��A�ibi�!M�29��$,Q9c1�P0m+b��D�}{cx�'�;Ś����l�LN��ի��.���S'H4�V@�Z @/ X��QQ¸āʖ����I'�>K�q�R�>�&vj����1�m:�0��y�vD�TN��∰.������=%�,� �8�!�IÌ��vF�_��#�=�H�l1N�����[j�/������iWdb5S����:	��lȕ��A�^C�P�<���ijaniiG"is��∓�6����������MI�4QF�T���v?�b��6��c'f]ΩwS�@�T�G�0���3fl�ڙ�03疔���κR���\Y�$�<7�dm�%5��z��2gj�޲�I�� 1>�MZyi+dd�=�8���`�nG�s/�N�̌�Ma��s���	��D��/��W��-)#P��(i}1-B�-2"˗��5$B��8�T�Ԥ��ֵv1W#:�а4҂N��b��$��shWX��w���Ĕ��
��,ķO�wa�p�Z��!S�Å�O��2�"efN]]l�~8�Lh-���U��g��v��zZ�ZJ����6�$�P��&�b],]�~))A<Z�g!ʒ	Ƣ;���e8��aO��2M.Bg�a,"72�ӷ�wj��E;S�!;9����)�Ŕ����zV���Ăk��5�ؖ�lK͙[���u��&��.�F9��0e~������L�x��J�� ��j������۶�!��d���ekH �}�GPk��˔-��L;99�޹Ė�ı��mA�\2��`=�� �RW+)H�XJ�\�J�hx�b�t^F����I�����q��3h<�b��%�<@+�9-��lL�z�i/�@d)�l��I�\����I9�Fi� 5��I$�B�Ԉ�gIs�69oiԼ�E���⯈x<4$)�%Z��t;Վ�r��n��o#EV�P��vK�Ұ�d�)3�i>��L�AYBό��I(ߍ�:N=��@7�H��$I{���:�����:��#�'�a��hcK'�:e{[)�,}/o�k�ם-���h�(Zk;-�j]3d��@6�f�i�e����JK�@�dD;xY�|y�Hbνs�L�����bfɕ��%�b%��̗i��$s>���L�a�Bs�K)T��ߙ�������,�gI}kVό"�u�F,ʌy�,�Xi�?3f�D���1��{���F�M�m�-T�H�tcK�0Yf�!��$R��$��$`W�t���12};�E���1f�!*}��c�V��.�LF�8�����Ҵ��6�ҤH�E��S2��z^�K==�Fh%1"�3�}����痥BK�F,���f�%˼M�d˧$m�:D���ڒ'z�Q�|�&YeF�>Q������&zMS�L>�5g�i�$s�i=�L�v��Z������"!c��P����?Q� �r[;�2T=C�s�3�)�_%mrx<�u�&�V�t8s�r���\�ߊ3X�{R��Pro��i�V�[�H#�x?��^x�y�.-�
u{CC�H��U���g��&j�7���4H��%�?Ϧy���hQJ��&���<p�A[}��ǔ�C_�X���\���ˁg�Vm@�XBg���`vD�})b�	��~��)�N2�yD�P�^*�'�Q��J�4[ �)ḙ0�6�2uʎ6%�W�4��>)t�qB���ĝ�t}�ܧ��c8rt�[�g��A��r�j�wd�Q8��T�؎��)�O��P,E�\#R�rr�jӌh9a��#�ˬ�J *�EQ�m[�rE�9�v�f�"S�}��6m�V/@����m�e���&#�i����<���Lz`��T��A���y��n��;7î��-ʨZu�)oAZV�qհ�t��� ��HXMj��Ne��2����9��L@Ԩ �d&�q�q��F��<�i9���F3U�_�dZ�̓<�"��,�`��������D�>F��-���RX�a�ZNJ�q"6m�΂ȔP�rjG�sI�C�mA�)X��}���Y�jUlԱ��Q�֚H [���v�J�x���BI���ÂdUϪ�TZY=SB�z�;��(���H���MKk��G"���־sK�-��$X��Ё�Z���K�/�l�f�iWm���:c����>d{�͆�2AJ��CP|W���s]f�:rT�5�g�:�ڶ��$��!��p[�^�`V/�2k���Ik���F $:����d+JOJk�ξi3�Ԓ�d�I�����2��X�:�!GyK1W�s��sLV���5�V�7k�5C�l��=W��G��c�F��v}�ڵ�Ej𭠱�A��5��4�e�z�b
 �Y�K�/-���=�K�w=�A�V"3M2�^2���r�Q����z��$ޟ���a�>a���JeY�\C�%�7�Ǝ��l��:�� ǔ��iq`e���2R��Y�N�ѿDқ��t�'�k��/Ą0��qO2���4Ÿ��酦8;PX��s�	ғa��P�h�x���$������Q�'f`��0���H3$���U�@�t�E�����m�:��M7�y� �q�3N�I�u8�t[\��k��)7Aj̀2���3��,Y��Jy���bmOC����=9���Ƀ���~L ��L��ҽ�B�T	��R�0σD���"X-�<��@�U��Y����h_x�?�c���ӭ�&�T�/�=��%�gk���=$��2�SDTQ��~"�$�R;�\T ��7|���"��=�%j�V�"�R��eϽ`���RJ�g��zr�{�g#$d�(w5��V��^�%i5F��j�B/��J��ͨA AɌ��~G&8�0�9�����ʳ�y�֦�$�L��D����ea�V�	*U�М��t�Z1��G�I&� ��(�*ᐸBU�TJd�fU��Й_���E��E{9����|p���ؼ�TY/��baqu���e�QY*dz�=P�W� ��Հb�ڃާ���ԱH�<d�x��oFh���D���U��N]����K��]X�L2������_�e?���:UB����6שW�~�'��L
=��$Lj,B�W��"�^�������;Mˀ��F�c�������x���P����\�b.R�=�C��f�ZMs,8�������5N��઺�G=�����`�P*�E���eP�Bͯ�c8
^��q�fʠΦ�+,���z{=c��!�G�F��N���i��t$u��B��(�~vm�t*H�I�{XsFF����[�����0V퇙{'��#��=1]���BwYN92y��P�w�Yx�Α9/����>�qV���tpl򒇏�B�lRTձf)�7�p5m)�"������գl�8ͣSp�0Zè�X�r�q��\��>��C��6��O��C�4Hp�|5����{�)p2�p��a�:�v�+�_�AT�y��OMT�d��F�A��
Za�� �w�����<��_x�/*S�����w�:{ѷӀf�ȉ��Ë/y�c��B۳�B&lD?s �w�������+k�X�z���׿x�UW]#ف�=xd�|/�?T����f�H�-*�&���������{-�nz���5��ort�P;��].C_f������Rϑ����n��E4=�Y�t:�."#�LAy������F�j�uߺŻ�6���)�L�I@�ATk��Ks6?%;������~q��M��zͿ�����_��W~$2�z�/�x-ݖM��EϮ�Ł���Mp��ykWz�l�S��_�F��n�)��G>���_s|b�-&jSqQ_��HNe0��<R��vr��_�n����6��;ܕ}�j��5�#Sf����CE�Ukh���ެ+3G.������OB35B�iL)i��"�k@�}�u���M�!�[��Q���d�3��cs^ ��W��?~�o�__��|�Q�>��?������؟^�'���H��g~��0$�p�+�����`o���s��ֱix��=��1ؿo�3�\q����*"9�/=�E�mLA�A8`�a��5�o�y��GF�?Tz�X-:�<��`�]מŠ����ua�7"!�+B�.�:�Y�r�k{Q��6��F��w�|�����̩SI�����X�/J&��5(�
�q�H5�-����Ё�|�&�뮻|�ٶ�m��f=	3��Ǉ!�������T�kZ��ԡ�;���*v����Aej�M	����s�LiSC4����<	�Ii�����0� ^9�<늦���땟�ɵ^=��7��/��e��Ri���0���C�"h�?���WF��sBd����{	^���!�;�B��v>��puf�4�k�����c|z��UW��5�>sۖ���yh�6�E�������u�w4�F�=���E����l>x����]l�N9�}�~x�͏n�d�U�x��O|��}g�|�����x��>���������`i�����Y�v�M�����s�U?�`!xa�ZC�]��Z��~������wʏzK��⹎�lB�g
�\ȝw6j�t0�PGB��J��-0_u�pDjS�v<4�����\3���_�ԗ��s6B�Z�_z�Ɯ�p�]Ĕux��{;��,H�S�tX>�a:?�����M�^�mx'���[�:�9�/���*��I�^�H��}z�.��'�
����{�G�C�����޿U�Y�m۶u�mx�U k_x�ɍ8�!O�)���:�&�i?�-*0D�|�~�;a�;�#_�߱&k��/<��ڭc =Cn����+�?���ޯ�M-���Y�?����q�����ಭEoK�y�|_|�Ω_���0�z�"`�\筸�,rf�%vh.�tma�����=�ښ۷o�3Qry�����{����{b.��B�ʅRU�(=a��"C�&EN�di��_ٞ���`���t(��^v�d�prR�����Y'���7 {����ro>���C�J#��y����<$�O��Q��C�݋��D�l�?OA'Z��D��ځ��ƴ�Ri8P`���G�W�1t�P�N����d����7��Q����������������P~�e�6|`�^��9 a�'��>u͐�����q`rq3��/��rJ���A�ˏ=Ƨ+P�E�VX�fk���*:��l����,��������/������W���ӄ@����P�4 h"$F�оɌ�Q͵�.���
�l��"����Iȍ�������W�	���#�>_�O�9��֒�w̽p�)��yіy׺]�X���+OK=�s�O����R�?CNC9��0d�'�,��Ŷg?QM��(�������.��IF?Q�1Y��IuRN� <�>�[-8��=��0��O�[��S���R�'� �H��*�5���e�'    IEND�B`�PK
      RZ	��} } /   images/bbfae99c-8036-4c5e-89fd-a87441410720.png�PNG

   IHDR  �  �   ��ߊ   gAMA  ���a    cHRM  z&  ��  �   ��  u0  �`  :�  p��Q<   bKGD      �C�   	pHYs     ��   tIME�#Պ�  � IDATx���{�m[���Ƙs����8��GսU���袍�i�4��A�("�q�6'9�Dq��E�HEVd��HX�d���&�Н��g=��n�}����ךs��?Ɯs����{����f�J������k�5�x��p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8��}�𵂪 ʳwQʄRZ����k��{�Lǁ�%O�h	*T�J�`011@��#�QD
*B)�@ FI�"4"L�Db4��L[�>T	
4AU0����11��*��J���N�L� ��m��l@�(`\m.@aW��7W�G�|������%���<�Ç?���p8��h��@K�J���s�H��K���EFi��_j��R�kh�,A	P@	`   �jQb���!f(PA�U{�B8��W? � �FE}E��z�T�0b��P�t�>��1�yPr�P)[��7���I�����>P�+��T�hT ��ۻL���J��ui� ��5%Nd?#��z�vH
U�w�[��}��rV)R�""�%' ��f�v�U!�bs�!lJ���x�/.��Σ�~�S�����G����7 xD������%b~�]  A�=��~l�,!	"bz���
�*�E �
$S�
t�Nb�Z�L�WaEM����DՀ�Ĭ
�h�AU���!7�(���?��˯���1(��a��%�۽�����]���$���}i8���U�5�ժ��T�[T�GE�C-�J��eC�����	d�VE�RM��F���dQ�liO~M�?'0�w^d^�b�Op�x<��L�$����3x� T"��q���/@%B���w���w��ڄ����k��3o������k�q����:Eӯӳ� e�n|�Z��	U�M"�7h�Yr��((W���� D��@U�����y��䟽��� �6� ���X��D%"H�T�(�R��0+���	|KLO�x��8L����m.��>��m.@aa�]�%����P��/  �Sm/�J��eM�7h.�SD��J�$_+t�RM��
 ن^X�f��@�aJ��QS�t��k��纽o>c8y�l�BqĻx<������{MH��sF����J�v�������U�v�+��K�������]^\��^��������ԟ��|�^�/�-�p����; t�0�>]=����_.���FD�[%���P�)	R
b�K)PUÀq� ̦���2���_�+t�;������2{��W�~N�D�DF���k��q( �fB8�g���90��2�d�����q��o}a�X	�@�>�G�ᗍ�VU����n�./��'�����/%�n���Z�K*%��Pɦ�T d�ά��H��Du�Z�9��yeӕ�����}N�]�v�W-�~��;?��c|���	s)(���QJA�fB�C`036�`6q��F��,��j�@�.�q�}�_o��v�y�~���g��W~Ƌ��Ǉ��q�`ڿ�_�o~��-������<�Β�o�o��V�|����D2��\!���!F\]_#�(Q�W�Y7ƽ˧3]oqǕ�\`S���"ZM"�� J�jTM1+���y����M`��P���ϙ�gƟ��~�Ke�q�1^\!��1��,���;�������/b�]�����U��HI�Z2 ��"	���`^yۨ�j���l&��mH:��@��l�
^P]���u�{	@��9��s��{<��s�7��.���L@��i��%c��؍6���1b�<b�#��E�0�+l����U�_�������b|�_n���7^^���, "���~����g~�G_�2��W����O�����%�v��7�i��|8n��[���R@*��PJC��`�!9���E��^z�U쮯�(��RU����� p� )�z�5���5ki_2����&�5���5�Ye.1WEO�����9
�'����e~������3������1ݾ��}�������o����!����?��9�.��T��9���I�"')�
�慢�B{�g�Z{�^IU��mt�Y�8��ieٮ����$��qԮ�0Q���.~a�9|*���ÌL���9�((#cF�P��BDĆFly����.�<`Ѐ�p��Kx��|}��[����/�~���T�O@)������W�������~�ǿ��y��/a�yʘ��b�]���o�Ͼ��2r�~��p��3,����4�P) ./v�$ bLsƓ�^z��x�ʫ��
� "���ӅA<�t����<���])U��kH��Wy��P��]��� �r��G��C�U�/J?�!�(��#���,o�M���#���#��p}�����u�П���|�G�|���������e��_�|+��*�Z��BHU��(t�ͧg}	yK���*3
�U](y%@hM߯��@���a�y��`��s����N_�8�@IAA���`F �!�b�
��1�6<"P t�J@���p�勏��W�`xTv���8?I<��ƿ�H���4��.��C   �7��+��4�i�p�x�xx<D
�:�ߖ�߭i��A��8o���� � �3��Md�H���#��9g�./����g�N	�^~��������Č@=Q�z�I��;:_���LV6�^�l��H���_׾6	�<vQ q�P��@���Y���q�� �o�D7x�c����@�P���/�*��A_�����폐����_�^�����Ayz�� � �J�h�V���c��S�w�Vν~I5!�)t�j�/%]š� 뤸��P���x=@B"��%Ct��@Q2��j�H1�Z��JI#2fd8!% `@�� 	!d��������F��:��?����R/�t�{C�o���6=~��v��o�~�qw����AU�RP��Bd�p�:s)�ó�?V4��9�ߍi���p��·m)�I��{H:@JB �%�'H�(iF>�Q�H4(�>�@cA�	�M7�i��;()D �%oz����q�9t�:W�dg�o�;��#����u��I�%�X�a���|����(�߮y�#!���@o}���8~vs���[_�N
��~$�}�y��޲,� �Q*��9�%��kXӀ2A҄��4�z�P���oYY����aJ�E�*��j_�*�cYXk�PN��l-(/4;��.�S*7����S�����	��IZ
� H�H�.� K-��"
5�d0�6؅+\�x�W.���xix	�0"`Ѡa��4���g���e��2���x��p����-!����n��K�u����9��3 �����͗���o�*2��O�\~_��o���O�i��N��y"�3Ho�Z 2!�#JN`"��9!��r�0�nn )!��8D��r��E@q���5~�۰���FFV3#R0Yc���Q�.DW��ޛĉ�~��P3	j��6��*s{ͪ���O�u�y�T�����UM�0(�X
�'a:��C�i�ݏ�{|����Ȓp������/	_W��/}�!l>���(�Z��-��D'@Dg�(D$��I�\��%�-h�Ӿ_|�U�v7Zy��1o��B������״}��;��"�ܴMȋ�iT�b B$�j�,�JBT�[J�A�X���B� �غ �H ��`@)B�6(��3o��4��4 �	�kL�c�O��g���8�0��s�Ͱ�~i������w1lw��t-����@��m�$�9���M<|囯5��۫W?6�~�j���K���U��n�O!�-�dYfhI�r��-E��	I,^.9!oq�y
��0n�u����3�4�c��ͣ�-bܘ�#��a�K�J��J�S���$�U�ng9��޳�R_T�9�h�EƂ�@�����OՒ�J�I9D����)㯕0��D�ߺ�<�����~������������O|�ʬ����O�ւ�Z��!�㿡e�(�)G�r�j2[���T�<s��qن�R�T;�Ψ*t���F��9��z�Z&'銢jT�4*���-���9��ւ�Y�]D@PD
�H%�&����Q�VC��H*�b�#Ka�]"�Lϰ��pF��~ʀ(
�y�&��M��7s���Y���t��1�� ~!����g_�t�3�C ¸�Ї��43�3���/�ٳ=��
WWeh���u0����#��̀�rP@b-}�j%A���BH�L@mX����D���Iָ���Z�X�K���jZ����1�}��p�b��`@IJ�A��AT0� Ί�2f�vD���q����Q��0E�t�c���
����v���}����;�y�%��j`���A����o��I_�"��>z=ݾ��*�E�'E��Z�5D8���h�C��	�@��|DIGS� H.ȹ@0�	ДQ�#�t � C���05���uw��"_? �&[T$K||�7�ӄ@������u�{��KoΏ9\����%/D��=����f_tN��;EJ�֛R7J_#�@uF)�e��{�O�����~����~�w~�w�����V���u��o��|���W�|��K�H���"G�L�2�lJ�%ͫn��1F��Ϊ
��w�yL��M����E)��z�ž6^O�:��׾�aU �Z"@�lB��;��,O�@����z!�$(J��ށ ���l���p0R�Ť���3bQ\L��-�����A� ��RB�v������5���������3S��8��"z�oso!�o�?�O?���q(1��%��f�tv"�w��T�Բk�a � J�s�a�q���	L#�iF�G�M3�:Z2r���<�������}��ʟ���G�q���D��2LE��FG�b�c`��B���L��	, )�M��`bb��Y��I ��H�tr��7�>½�
�����_R�U�Fji����P��
U"����V!�K��R]
E� n�b#��:�Ah�t�����p!P �����^������ 8>y��h
n�S� xh+�Q
�60C�~a�.�J�s�JB��g�o��}�f�g��]4b��� )�����/�9^
�Hy@�!��H�q���7��oW�߂r|]U^*%_�f�P�W�Vb�%��@�y�e>"�(ǣy���-e���'@b��%c:� D�4�e����!�@nn��gL9B9X)Z) ��oN��%�T��G�ÛR&��!��Xe�$��nғ�A+��.R�m�e���Ξ-�K��%�i3 c)lT�D@��H��)�''�o.����nz���O��#���a_+|���f-�a�0o����5_)�R�Ũ'�H-+SA˃T]�oQ�a���g�8M�X�jU�X�6ֹ-���s��2�kѩ
Z)�wR��G�؅["D�Ь(�0A� 6A�(g(B��g��#B�dU*`Q����)^C�
�hA��43��A�!��A�^�^"���{�BxF����D�%����ox� �q����ՌF��� r�0��N����N3�W��z���y `_��"����.
D>����d�"ø9��IidC�qP�AJ� �1�C��n�	1��R؍X�S�4A ��(TsE��*7�\5s���C��L꒮oZP�7�7T�/IAbJ]�i*UΩ�Y�(DETUE��Q��q��THJ	�E��,Y@9�EU���PJ�&*��"���T�\��-�˂�-Ƃq,�~�_�9�B�R����٫Z��*���l��r�^�3=��C�<�������`�hH�޽P�E�#��HyՇy��\i�;���9�ΐ־Y�'ת
J� �(%[-�<��#��M	�fS�R ()4%d�ӌ4O��0#猔R�P#�b�R��0����f�� sg8툩9�M�5[���Kύ& ���K�{}��$ԭ����ԍ�ƪ��ηváv�_=]��p�b� �d�I�oU%��w�VDE�n��2��ܼ�i\����zV��*�ӻ�'{�q�M���/i�sH�G(gh��V�V2���>���@��L�QSƴl�N�t^~��۷}JQ{]/1��Q�&�v���^N� ���M^[�f��FR�`l8��#v�E�2CHl�Q��I�d���I�zp�`��DDe	 &&��Tn��u�b@s���\KE2�L��  03�Ja$#��� V�P�C��8&���(4�(QS&��L���U���(I��+���� ����k����v
�<;��T�i�����a���2���(��r�BsR��H�L��HDL̡*_��i`Bd!��͆i�/]1^}i
�U�K��q�u�V�����û��|Խ�6L+MD$���Ｔ}L_՚����R/n�7o+%Y6qVe) e0���([�DDC9BDTPP�([P�P	[`���P���VG��"�%�HI��R��Ǵ���V�!T�T�c֜7�������Z�̌�{5Z�v<UHUI�����V��b��*K� RX�0����b^}�P�*��g��S�Ħ�i�q	e>�oQ��d�Ϥ-�Rl��������
���cJ8���%��ْ�b b4�:M{H� �S�-iM�@cS���YS���3=]<4e�L��&��7��D]Q�2<f-��w�n.�~��G5�,"�mb%S� ����Cx5���k���n��4r�x��O��Z����~��C\~��雟�m�������'PI֛Xg@��=��F"�j��V��w~" O��~M��S4����z�}�,���歯�f͆��ڇ�d��fc5/{TƆ��BϬPeX�2��Q�D��p���� +#h@�!����!?E. �ƂѕD���huRTC��� �"�z��`G�� ��o�����Z�&�Qz�w��y��CUf�<eL���O�xrTd,�X2B����$b�:
�xf�<�3{�D*}K1�ĀAB���0!h��̀a�������D!�����жt����M޻��o�[}����F�,��'����ͻć��ď*A���Rt�-^V��$��%b�p��[HA<a�`� ���tܢ�K��щ�P��-!l*1AF��lbM����l�=Y���
{?�x�=Y��k�
h1o��Ĭυ4�C(�"E���T{OT�ԩf])tj��u{#I���|����) �֬�~��j��|D"R��<�8���8D���M�l"B$��ʼ� ��7S�(�i>�϶լ^�n�ﲹ�l]���{��*���F��* �:�et�볰<+2O�b芚���ĕ(�Q	Py���P��}������ȳ�O��)<x�[�aǇV��~����@���4���n��*�
��5Ͻy�B���4��*���{����z73׍ghq������K������������E1[���
2�P��  ���
��b,�F:� E�Rz�A+0p(��\`��y
(]Yk5����C#��jV��!�׃V�q���#�g*w�ξ(�/pW�j���1�$I @�3n�7�`�@����D�;WDP�@T0�	%[�b)&l+8�b76RT�	��U�h�\�	~'��}����N�25�6��~��	Z�"�	"]��l�
�{��)T��!@��t��i��#Xf��`�
@cy��4@C��-hs�v�n�p�{_�U=4�¼(��8�2�M�[S�XN?�m�(s�5	x.�5>�3��j�I�z�K���O�,=f�{���'��=@5�\�]q�P�#����JNV]R�0��V�V�3BP�t�����^_B&3��R�t ������ߢ��h��t%��2�O����T��^/�k �Tma��0�����?{�J�KM�CϷ��r�若�E�� ������������'���{�	�|�Sx��oy�g���R��޾�gሇ�UM���K:��G�̖"�f�Ve^�~	��!7�l�n[��%�ӂ�-J����ן�)z�+��O7�J�wLZ{Rj���5�X���ʜ �2�H
��N
S�\@�M�Aњ�7Ȥ"(�}ge5�t�@��r�1�A��`�8T��湒V:��}�*�%j�ΐ�E���m�"H���:��`�ύjڽ���D[̀�� �#O�,RD�l1gV�@��5r.�sF))���!R�e�0�-."a`���UjhדX�3���=(*x>V���-LY��u�� ��=�u4� pT&�NвM7
SX��0���vL3(O�<�'j���J�TD  <��:o �%�`�ov ���^rZ�U��Ր�5-mMZ�ЪL�p��Mq��g�n��[Bz��֥��m�h͏��_H}F�Xy�-��׽�O�}��)��a��$	��L77fP��
�����mă�s��2w�v�n��Q&���	6�U�!��o�N�Jj�u5��]�r���5[��ht�ʘj\���AlD���^�Q�2�~�*��~`�L3�j�Q���`���69W`{��$
�����O�G�+����`��e|X�S�
���ޔ|�'$�T�<hIF�kF��PG��r�V�V�̓v.+ֶ�Im���'V���wS�k�ܳ[�u�z�<��/[�]ey�)��ԪI�l���w&�v�@m��d0g(�*��%����6�%P�Q����4`�r�$3����л���ٵ��^&*�W�*ШUi��P�,lM�����Oj��w��(W�kJc�͆ ���Cf�"(U�81B��� �\��{�V0P�Zl��-×a��|Ļ���u��
H��O��T�C��]�rQ�͋�=����v��(��b�.�`���.��9�ƺrD��L��Ϫ	(
� �	�� %�����T "0,��T�2�)��!� V�._�� ���M�	b��GX6�+��:ٻ��5m�*��Z7�6���S�|��β(������h�Z={ċqQ=z�RKK�2��,Dl}�I��,N���9�!0(0r��b��#f�-V"I���`I��7�f���ۍ�<�?`:$�3dN����z��
�:٫��{�����5��x�M�wơ1w"+�[��`�G�����\�3���}4̌��OU�#֌�z�a	J�������9=���G���'�����q��gq�!m@�S�7��T���%����%�XӒ�e��l-=�]����+���f�����j��$��Ic�٬R:�컀&+D�F�¼��,����*�C5Fd@i�DA����2�b�'�f5+�Փ-( R$�FիoP��(2�5��Q��/#c/��2n�G�A���vo����Rf�;2\@� ���l�r�@�Ӣś����O�\ʲ2wj���k=1�B�l@R0b�u��	9<�f(P�le�2Z�p$F(&���d����Lur�Ֆ�R��
�12�����x0(X'�&�-���.���[����J	P�o�Jm�tU�띪�ꋵQz��-g�R�N_Dd���	:�V#���Wg��
��`L�,IrU�TD���*
���n!�-�b��PF 5�����B���O#�-�e	^�@lFT���<'�6N�5׵Z�ֈ��贌����3�L�Z�ZmHͣ�&�+����o�
o��vT((�e!OG�)a�8B�`�7�W�����O�<��֔��|�s�LG��"6q�V�K����YyY�nJ����^��:��*p���T���85�~�4�3�<�ET_������J *5�*˥�v3���k�$9�/!��O����ç�K/�>T
}z�H��'�|�Ki>|���:!�)	��lJڒF�4�Tzh���Bk1�"[�R��tE�uO��V+�����oS�M6,}�[}d}��x��
��!PH=�k%�����(��`�)�X��>6�	!��MHP��D	3� �z�,G� ݮ����,c�f-�|q�5�u*���m�cB��5���+/H� �������Ѽ��x-$R�9�T���9�Br�� 8��ԗ	`A���
)3�
���2z��@�R���RlT-�R0� S��`?r��y�]>�k���ݵߴ=q�e6�Z���<�~��{j��mˡV���Ȧ�+���6*����D���̥� %�L�3�c�j�V��?GS�f`�	 {!*��C@k¤�A��^I2&��0)jߘ�%le�w2�K�C<�<볳ؿ���[;�K<[����V���.��*!��m+��Y0�*aD
D[WHE)���h��!"�3?~�9M�\I�a`!������./���/DH�1����iF�%3�焠-n^�U(��Da��O7_Ջ���׶6'������ڴ��pL��idJ��.o��oK�]�����M��`�Ř��>��9zB� ��o�7_��v����[��/�>����Q誊��/!�Ã��͟+����<�J2�\l�o+�`�D¢Z�E� 5~��$�d�F�-�k�}+v]�D7VX2�W^�J�T����i{�	�槣�!U2�bk��Z'��`�[v��kw�~�%2� n�>�{�8ҌIf$(PM�#�f0pD�4� &�����܎$t��Q^)iՓ�5������Z�t�i�a=�R�P.��	�2$)����<!���JѶ��1FcD@�hID)�T��"P��{�Rޥ*-�K�=�z������(�^�VN��BJ�F�<�u��'5�AD�O���[�q[y{FEP������PB������ws�fԁ��B$���0K56YH� P��8��1�8�ᵕAB�~i��s^���^'���w��DO�ZU��_�.��B^����!��?tf�����0*~=DJ%�>���Ŝ��[�yBN	77Oq�&�֫���k��/�q��BDPR��`���'����'8�(s��4M� ��j�����@M�yW������BS��o���3�(���Bn����\������nșaѪs �_Z��%�ތ\�1�������O��;�����]|v�o5�&|(����������9������<�ђ[R�1b��%�Y\1KY-~�g�7ũ?���@��y��Q�%�ף�(zvh���3!��n�;�@�����7b�線�F���J�Lv�"@z�0{�v@Ĕe��$�P�g5�V"w(3&9b�	%�`W�}��j�����#@JFN�QJ�`��P��r �լ����h�"�(�F�׷�>k��F��Z%�2 �)f��~5\��@�i&���y�R�#�1 F�u����"�!�keA�sQ�T�Ů?FFL� �ϧ�q'˵�H盡��]��8`�ce���4�e��1&K�9��
϶΀e��ʘ��a�:im�|ʼP�T��R7��{U�x ��h� T�ʆ�5T�/D@f�<IP	�o�������c)��%~�i�n�/K��C��nG�V`(j������k�gM�=�S���I�Z:o�v�TK�<"BQ��������equ��d�>}�y*H�#R�8�v�ǓgO��l0������)%��<�\
�	����Gf��%l���7u�,,�%�ô$�َ'9K�@�r����:�җ�3Q��6�h5Z�:;-����)z�LY�u�2]�r=� ��2�������Q��|y���ǃ�+>,����"����]|�o��S����<}ea6��՚��I
�-~���Xr1�doz~d�z���������j-a�3�W��X��L�L��1*#��e���5_]p��aM�5�A{G&�L`����Q2a�#2f�Z
 B�� ;$��5�02�x��F��x����0F�U����W��r�%	���,KZ�v���߮�sk�c	�F�.��j��S�-	�Z7S��pn}�T�JAI�s.AB�H� �(IPf+�4`�ڎA�%F����m��J�5o�HWR��{�'�����e�`�t��S^�g���JʟP��fL'��d��`��ք�Z��e��["�P5LXZ�F��s�X�n{E������9ke+��u�v�1��Q^+�sZ:A��.9�gJ�mW��E�����]��wj���/	5����p���J�Q����R�tx�iNl//��G^�~������ FJO�1��r��a�ʌ�xDJ	Zex�)�sO}���a]���㥯�k�;"��Ȩ��\^c��V��$����z�S�W����I�z�^#3$��6B���?���/������}��O��cߌ>p��������7�v�돤��?U���J:�%�D!ɐ�{2��R��s��r�~��K&o#�j�2 �z-6Ӕ���9x�ڼ�x�h���z�,����|�r-be(b����q,��2n�P��0}��S��j�6���%aFƬ3�L�2c���l�!�pG�C�ц�l ��xF�R���,�z!��OX])t�$����x�,�{_�V��1w�J�
��� �1a@ҌP
B�Z��X )c.Y3rJ��>�gD�F���E)+R*`hQ�ڞ�4�*������S_���5��[h�y��������0+����e"��Q�EiA��iz�7&2Mlg�$��0��T#+t���Ĭ-�ь 5�Ό.!K�5�l�n.�����ڪ�_)�x�ٛAsj ��v��
���F��I�7���W�S_��("]�o���9\Փ�����QE�d�C q@*�<g�R.8'l6#�FpQ�qy}��|�u���x�����}�� �i�8L38D[����	i^�,����3��s���Qp�F��$c���oxnI���J�\�{j5�:+��8n=1L�����\�e ��L	N��
I>�����0=}��}o���x�o��T���%���ax���(��G�|T&�Z��6�	4Z��K?�Lړ��k��S�Qd�� K���Xka���Xv�2?��Kq��/8��V�t��=ʿ%C�6��"F���������ѫޓ�:oAT�X�M��Fւ$3�L]�[�j��z�bε�e�vW���8>@���:C9#�Yp�����S6���εRWt��}�L��n��lb1�w `�)،f�
��֖��c{(KY�KR��X�%�eA��`�C�hQxUkKlԟ�n�?m��
��;Վr���G-�g�hԽ�h�*���! %,^��>FcQ�GҌ[��5-�7�޲��%���q�8�&�ڡ�@�Pڹm
�Ң���[(Gc+Dj��T���E�:/����K�����װ��Y{R�H���3��(��#pzx{�W���2o�C7ԛ���3*�[�@ss@�qq�4g\]]���#���8N3�d#T_{�%�~�d)x��cd���T0�qs{���{�a
��rFN�ĠYd��lRks��t���8Y�;����K���:�������H#���ۺ�I�Z���~���B[�f	�"��A(vn�:m?rI b��t�^��/��>���;�>��ۿ|`
]U������_���{~����h>��2A$�g#����	�j<]!@� �Z��&&�-�D;�5i:��d�V�D�P������e��k���y�H�b:������;�[Љ
;�Ӈ:�KA1��0b[�Q��)����ژT�@�2*�n�aP����lY�(�R$HP䈩�"˄P�B	�C�Ad��$A�%=����!�xe�j�!<d�Bt���&a�1)���u��{+���E��qq���ŦTJ�BEj��"�pE�����焒	4bX:X��Ա�@$BΊTj�
� I	b`��`?�΄cV0�d=�j��P�h�0�e:��I��v% +ͣ�̖��R
��.���?ۗllPh	�U�	`LK)(Z :!ȡ6	1!�4����$"����JMk_]�F&k-j]�
��l����������4�����	����E�֑ �)YIT��ֹ'���ւ����v�m[v�,�Ѣc"]�-L�:�gevF~�>5�n�Y��+;��i�����w�l/����ݣ+l6�4�����f��^������	�b��<���,'�x8����r�m�{5M���#'
�}y���vΔ�q����L���g'���t9 �o�u]����C뫯'��Z~�U�؜�j�$��I~�������������߂����|�o�-�������=���I���t� 5���,Ѥ��-q2B�Y�u�A��ن�W]j��.�`��O(������W5��w�Z���|�$윾�Y��\� ���7}A���[�U-.W։)�M�b���,����f9X'�b���-CY��?:���@��:C���L��E��������� $�Z�o����,ٺ
�nNUa��ߝ%�����D�c�E���m$"d�q��fQ2�T�p HY�&�D"D��`���5z*�\�X7-����o=S<>�K대dzZ�*ζ:XNH�ԖF��=��c��Z9���a��\�Jw�)Ag��^"E! J1_�,fK����rWB����Lw��(�Evk76Hm?��[	(��a����e�`�|v�������a�Ӄ�&�E�5�Q��f��J. �}�j� h�H�S�f8�Q��q����z�-sga�Z�jkKZR��i\ (6�t6`ETPJF�'����#����a�-B���RJ��v��	2�9c�#a�ݠd`;��n�SB��)8��)M�P%�J�!�,,sKe��{�x>I�<Y�;G�����z���c��3���Fw�c/_���>
����:�	l���a.�24-�D"�%A�d��_���y�}+�>�<.}>0�>=~��똏��W��GJ:��Ɇ���#���T�]J��Z��5�^��K�.ٱ���ߟv�[���`
y�1�f�)�=v}rg_��(],����p
�u� m�.�bD`
��jrגd�(�H�ſ�P���EfZj�U�u���Z�EY��U�	a�#�	*���H�,�ea������DKM�Z���0Е!Ж��0�H(�\=j�GV@R��j�s�&��J�zܘ�$"g˼�LP@����Aр���@V�����L���18��ߺ�qCN�����CS>��;���@Kz����q��ǵ�U ���mF�V�3C�2їw_�Gv^�a}�hM;��Ty���"���d"Y�Bɦ���-=y���=�P��� ��"+O�5�i}�W�\=c�)�O�w�V���*I֝�t�m?\��f1�g��i��[_��&@5A���^�j� ˄i>b�#�`�MeZ.���߁����A�f3"��'X�RPJ�dWǨRs�Ob�f��f��}u�V�ק�)�ޟ��q�峽�����Ým��xr�r"_t]]�Ƽ
 *���=.�2�1���O�g���?|�����	�������UzH4g�o�B��$�w�:9M{)Z������dP9��E���U��Xj?������[��7�*rfMU���ݤ����sZ�Z2%���0%�Ɇ���&�B7Nl���i$��5��דs��SR˜O��:#�D��#����<�;ͳ5��d�&�N�������`j�nBAd�z��^/�s�B*�lXw[k�o����[���L�o�m��a� �%�Υ�Bd����T���U��CR׮������x��w��?���Q�]� �����s��vJe�X������֙��������J�+b�!��i��[+�:e��#v-���K^Rm���/�ql�^�:U�
ъ�4/{CZ��v����7BNAulks�AK|v	�-�	�>9�X��*��_���-�R\
3n��|#����)��A�@ ������vLs�������^sr��@���%��n�#�<M�ӌ� ��<�w��u��{KM}ϟ�����-���'��:z�*���V�ja=TÔ5�Xȥ�L�Kӌ m��@Hy�.�����|��o���>�m��'�s5�Z��+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs����|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�f:���E�s�.�L����)������@��w��{n�<��D�^K6�md�c�pcs��yN���I]�$�����i�!�����9�x��=���b��ko@�[��E�S��y�a1�F�bf���W|��	�64졻V�#���޵_���d���є\[���0�h��9N�	���N�!�2�}���2c��?�ߝ��
���{��HI��z$��W}����7S��o=�|ֶ�����]b4�3R. f$ʠ̠\@egJ��%�Ȼ=�T�4�h��]�8T7�1�j�{ȷ#�i���f^���=�d�w=ܲ
	�1Hg�|_��O�Zb#��cE-cm����>AXj��T M�Z�iF��3ي{o�GE�z�E�8c�v�7�n�6��e��I-����#qs��F{J��w`f,�y+ �׽S��=Ӵ���Í�����WV��H7h�!�kO��6վT�#��N�l�N�E��O�2��e9~-�����!�xS�U�׾�19��?W��NH�w�ȥ�"��x{a�p����Zĺn���|r�j������!,}��}cu��o�2�T�6�;�n���1tKY�&�!{��1��]�}zߺ�F��t�*���ER;�H�t����ǯ����z��d�a��x��iW��Hcx��-`�*c�&�b�ns�z$�o�g�{/E$\#>����ЅQ��HIM����+$'�4AZ2O~� ��yM]#�ߌxn���%���L�ځ��ہ�̣��c @�b^�l��1.��cch��}=��&4��ƒD+oB�#��G=t�b��O�Jid�m������>uʫ��C��i�&�T+n%+n圁��){4���g�$��J��kB����ͥ��V�ƃ;�:�J]]w��{�X�?�:�&���=��������O�m�j���*V�����*C�=,�!���*č{��UD��������ݣ��q�=M�\���58.ɚw�iY{���tG����U�-��~���7�O�o~�e���� �il0�C��Ъ��m-r�� {�sB*;P�~�S���� ����x��:П}�{���9 ���r~+��H�X��ԭ4���}�o�@j�#]�^�*$ [KR+�#��W���s�Ƭqtݱ��m�|�6�]�ݲ$�|zYh[=�=��{zQ���f`�{CX��]cX=
�եz�e��i* 5�¾Ag"$����LDA}L����vA��!�Vo��t�2vۤ�o����j���ĭ>�s�����Jk��\,fqO:5+�Y@�����`�083L��&1���e0+r��guU(ߚ=�/��N(d1���WG�1!� �wX��̽���z�ͷ�kߓ�XQ�d�:x����I�H#W޽Y#)���:M̢���t�܈+�$K�d�f�]��D&I^�h9��� M٢>�w-���ugQ��������[�˼`�ŵ��ͫ��}{{���F?n����%��m�4����>��	�s귕��WHպt K���S����TPe��Ċ�#�ہ�Z3!g��tlW}k�Մ,�c��xh^Dp��Hy�Ϙ�)\ER-Z'	@�>Q�ڣ5↳�BU��?��7�������a����^{3D��m#�2ڂ\�������$"�w��;��9�8A�
��r��\ (�N`ڻQ[@y��Ȼ?��?�7�����?�7Ձ �����_�9,K��n�JOr��ip��0���P��NԚ�x!ء�:*K{���G�������c����_���pc����YĲ	k�Yi�L��M�0i�>�O7�77������ɼ,�l{H�7�Q�L�F&��5ܷ�R��0�> �c}����5�%��� 6���m8�/�Nv�j�$~	��A]<a�:s#\WEU=������hJ��-R��y�x>�Ɋ���p�4N���*�f�kǆ��q�'�:G˩E⑏��5�QJ��E��k;������0<�/tv�ֲ�"�PuHޓ��i�l�����'���f�71�:�^��)!!�Y�F�i��^��̮�X.���R�.��*VX^�6�Zl�^X��t�Ϭ�$C}r�n�I-��g�����]��^�W����X�����ӫ\k`�f
p̌R\��>�4�h�v�UR��5ۏjkX*0�Z{V6�͕dG� �_�{���P�u9�I��E���5r3��#�Q���-b7�"]���=j�Q�d��^6��SF*djp�<d�X�4y�������t����w�Agq�����~��K���7~���NzE~�HY���h2�7���rZ=��a�]�o�2�����,k���m�cV9�߬�'76Y�hm.pϫ��Pݶ*�o`�y>���r��e%�y�͐t%� �V�:B�6�I|��9#�y���@N	3^T}x��i; ų�ÓD����5�{�!�l��彘,�^$�)2Ī�uV�M�M� r[<�A�J��`��ŕK������J������@�N	�^��
4��Sww��3�^[/���ӄ=�8��I���Z�:�����������>+�X�����:�^�u[���՝t�+�48�b�/��	>�N���SO�)�&9�5�~h+e0'��m��R�C1��ٌͨ0���z��A��g�y��������@"t��q���z�7�\\��Ū��Vḧ́�ך�_l{�=�$�ު���j\�J���r7������f`8@�V�	)OÐ�V��d3�ن�����u]�P<m)^i,zlp]��v��{Iלޮ�n�l��gA�m+���Kߺt��"������ϻ<��2��	x% R�(�<�ly#�I=�)!BJ�א��s����2�^���A��xS� P���o{���?��~�����|K%��M~W�̓���0��F�Эƞ�j��e{�����@�l��l����]e<�}'H.[�19{xh�gW�z_���
�0�y1��؄�Z�W�ZG����f.���X7��X3#b҂ H�$s�x�i&{���3k��!^?K�ٔi��@���u���:�6a��#^6�x[�sU y�V`n ��y�P������h��=�f���\�b���m��	˲@!�rBNdS����̣*��|�K��]$�W�����f׍y�z�c�S&�������خ_���[���ӱ��f=�����}� aW��e1/�<$��{�잒��!�Ecm�׾�\���@+�2��<	��$���,�v_�쨧��K�6�MX�/����ֵ�][�_;����@�/k�}���~��x�ǟ��vcٌ�_����o�=K e��6�~Y��� MpCI��n͢�Sbp���^Y,(@"F���ڈ��LP�H �)��M�3�،G�{(6?\1�q[�G�H��U�p��9ҿ�h�����8�8��=j�w����!�c��E� W��8O�#�8'(gP��T�<�R�0=��~2��+ǫ{�=���Q�y����~��﨟�9�����Ͽ��?�����"G4,X����C���IA ��۵J�ԇ���R�^/���O�6w��鮘�mB�:�D-�	�.�V>�sQ�Jzh+���R�2]�!�ILloߋglZP?_��IU��b��EO*�����t �4r��mU�g�{}�ȉ�h۞���?��26�5f�!Cү
�MR�Q�Rd�3��n��{���K2V�,��V\^6<)�L��Vۨ�ruh�S �U�d�3 ���խg�!e3D̨i,:��յ���޻�cܧ�g���ՙ��z�F�9��SztC��9z����~���M�A ͞̳�1r�������WkU�|4e@���zw�}-[�;�-���}
��]�2�Ț 9����ģX�0���y�\�|���q�����#i��n?-g��=6�k=��n�z��X��kU���4��"�%'L�	9%;�`�L
挤�T9	@�l�Fk�4r��CY��
z���M�B܈�\�H٣~�������zQ�p��������7�����zU�Yn����n���zU���{�*m�ל���@��(Д�����7�\��mJ{ ����ɟh��}���aqޤ�it"�~����Ư��q�����OO	��1�H��֦�^A����e�B�aH����#T�k�]M���C�7��ƚ�G��.[WF�yzŪ=�ݳ{�_�(Z��Z�V��Y�_���'Q�VJ�D��Z����3�0��t�6v�����"����)ﯕ֜��ٕ�n�9n����X�g�W�ۡ�s�.w+�:Q�M��s���e��+\���-S�n�qy!x��@� R=�n��j/SL)#1#�Aa�2RS�g��L4[;���抔3���L�\@<�6����h��q2���zR�b���M�j�7����Gd���{�CZe�EٚK6.b�֘�(2sF��BW[ߍ�
2�L�T��y���!����sF+tqt�.��y��@/�Z��wz�Q<�]O���zM����Y@���U6��d�{�Q�p��l�x3 s:o�!o����{�Z��li��~�4M`2�k��b�dbO�JV1�'�ͧ�l�*���*cؑ�v9EWEi���O���Q5�e��`|@�����ݯ�*�D7��X�vO��,cF�f�z=Ł�ߏܻ/w.�^�z:]�L}w6c���{p��yO{����0s��e������ `�(~���ެ�it CB�s�(�|]./~��<x����0��ݽ�q�k7�M!��湨����z��u������X���æ�lv�&44���%��t�9��#��4<�ѿO�屛��L�������y�Խi �40��v��`$O(��K��;�m�%v��IM>��=3*(�9�++	�������ٟ{� �:Q�W�JU���QEէn	�������Z�
hJ�1-G\��oy�Ɗ��ZQ[C�L���PB.�zf��y����&X��V@����ē`i���PJ��eƝ�~���W��&�9�f�mk�p�)*�zlN{t	MҪ7��w�Ev������aHٌoej���v;�a�r�l:�P�6��&���N;H���A@*;�i�@��'s�tq	=��.�8����Ji�n��a3�'7�ӣo�`$�\9��#���l���#2�kH�+���p�ѝ��Þ+��I�^���}�Wd��[=���m���b��n����N>��B�x��-��V/n�����G�9m���\�\zAl�
jd����å�>i�H�!��G��,����U~�������H�)Rqs�~�	�ŏk�EG�f��;@��kDJ��C��Ɣ����2퐦�T&�r���i�������S�����7���M�M}�w����s�(>����������K*�	Q����˧���9���e�ՕP��=r`�ʔ,TBCAZ�^�Yվ S?�W�����z�h-�R�ԳC
O���Gچ�\�]�F�����Ⱦ �(�a��B��@�)���j���[�	9�0Q�!gܚv��.pQ�8�=&-��9!��vJ�>'�Z��ۃ��d�ѣ��MW�z���am�{# *r�P�̌&�|D�'���l��{��	g���A����V.�Z��ǓU�i��3�
�Q���a���	mO(��e^���b��dnD*NMq���'2���t+cAc=�t1��}3|��^�E���t�Ve�*���E�x��;��}^wJ}F��NH��9���=\��&{b��кN�y<�i�`KM`�ВВ��!*�߃�'!w��g0JbdΞN�ϚR�y�<��7d��(�ի����U�&��[����Nڣ?�Ag uY0��=?SA��K��郡l*[�N�
�� M7��6�<��#�,H�L�`ڡ���&�,�V�'IR�tEj{��p<][$*O�i�z��CS,�tid�r;��?�z�9���"M�������[Ov�)�S�Z��E�v��6y�.��3aҸX#�}��+Fl_�}��
'���#�����-��:X��D�+�?��2A��\,���`���:�>ޖk��G����S�7�o��C�3�0n������^~��9ܯi��+𣤺K������|�%՞�@nM{ۅ􇗺����V����V�@�W��X���K��m����xo9a��Dmآ�E���ƿ�W;���	9��5�o]�@2#%�BJ�����[�`���T�����3i�e������%v(v%SvO P����=����U��>%�BA���H�_o�̬Tv�DBDJ�oӴS����'䴳��4�ݑ[���Z��¢�V�dJzJl=����`�k(�C��&�s<����&03��Ќ�)�J.���-|�Kh�Q���D6��� �	�+�d��'2�'�����б�������Ƴ�j����ѾǤ;����/xލa߽)����?�+T��n#]6�\lP���*H:���(B"�5���R&P�x�M�4�����m*����S�˧�r@&'�V��o&���5ZU��`���Ƭ AM�A�H9�%e&eb]�E[�*M�*n����������N|�����M�D���'�UIDIUHd�Jċܴ��}��.��0�X�R�)_�̱��� ��?y;��3)Ӕ��_@�p�X�()�	cވ�Z_����dެx�@�!���RaKM�}��M$��IU��u5�!d�(�5�;F��(���F��7������7�S'=`�=#��h��SA�%���r�;�:��ns�3���j�������\��|Ͽ�����?1�2: ����_�ٟ��˸������{�=��$���酪���k��+���q�����f�KI���ja\/"���zC8b�=4z��r{@������G����xiKtE'�zPTm85A�#�d�c����>)I�"��gMH�(^�iyfFJJ9`��\pk���t�|�|@!k� '$0)Zv�>�����������S#JU�-��DG"����> ½�t���!�'�{<pՓ�^K[qF������
9��*�*�T�lҞiwU���v��}-�:�'ngpR�Xt�@p�GiIN��2��e�t\x8N[D��v�D�����E#B*��pk���-­���.����yL��X r��k�ivD�2���MWA���vf����^�E���Y�U@�!��. d*����
��Ҿ��4%�\4��!�"������3v���O@�L��K��'�O�佧��̤��&�ĩ1s#BUEm�.�<SJs���r:��� >NJ�>щ���隠G �rﵓ��"h'-j�,`���W��(���p��C�])�n�����>�|	�U=�&��-mr)��փjۋ�I[+R[��L��$���"�T��HZPX�XG�\���).��)��@�KL��Φ�ժh�J��Ac�>TB����H��nl,��&P����=� �
�V�Aɮ��;�ױH����}���I5��u�g���)#�؝��*S�g���X�H��{��}�E)�K��7��v~��,�Q���w�9���G?���
~���=�f��˷ԁ ������+��q���_hy����m���<1��k�/Q�"%ki�&Hb�0i�N�:���*&X�ܛ��x=��hxI8������V7�U�C&`l �U`Q�PSA&��V�'�W ~�0)R�P�ȔL�L2�0�f1QA��r��i�;�ܙ�`���<!���VA[`�ښ��Y����T���<�Ӄ������5f�� }�2^d�<����h͉+���ݾ*s��n���ҔX.�����2��r��Sʍ�y.Rk���&�eB]
8=U�߯����wcW���������T�E�ITx�j���P�'n)�4/x���Ǚ�JΦ���	9eH3)K&����S�>+n���pkG�mFW"D���+����}��6̨��m�.o�J]ꛣ�^�lm�Ex���~��Z�.���. �Z�����	uf�(�H�V��݄S�q:	��)���gԚ���%��ٕJ�n/|�����S��#_3�Cb<,�����_�į xE��,*ߨN/��[.��[ޕ�)7�,�rc��D¹4"m��kd�e�&Mx7)�De�k�,�jEz�Qr��m�@��r}dL�y*iJ�K�Xu�mn	@Zj˵�,�%�9Km���V淋���R���|�H}mym~B��Vkˡ-ׅuIB�mAʌ�����q��i�����B�N��]ɸ�`\��КE2
d)�vB����hb:]��HPP]Еۈ H��u�Ż+]�����dE�"����Q�;��'�#u�BDS�;oM�{爌Z�q&�a>�@0{�>���>xe�R�#O{�2]q�-�������������R�9�-x�v���Ox���_�{��Oѯ�ҿ���A^�E�� -&�)&<Cb櫶il��R����D��dZ��\���lz�{��f����!���&N��@2AQA3�넂v���z�����+de
��M�1MH�=�N9{�3�JW�c���].pw�w����z*C9!��Ҥ�,Dt��&ί���Μ��S�\N�O	��*��9O'N��ʇ%]ޞ?�3?]�|��r��R3���֟Ih�J���n(������-���Vlr�js�L��'���������9\\�5��Y�q}��YQ�KD�[k���i>��c��[A*Y/��P8=��J��e��yλ]�23@���5��ä�ĉh_wD�/3������?����²]KοNە�9���D�`P���F�1Е�[�pV(�GE�B��:V��� �MՆt:i�_B�	����Δ���K�Zv;�ۇ��R�I��x�s�j��P%���y��SO�r��xI�o�i�Uʻ_W�/���
PK�%���VJie�qj<q�����7e��[,�"��y+��v��	�fc�T2���tЗ#�X��'kgj3P��5�S�L�z���Pv�L��Ί4�EZ�5H���P����"�a������u��Xj�3Z�2�_��m^^���h�۲�g��nk�����T��z(:CeA[ԥ�-���e9��#)���.�*{Bk��:5��m� ���־�D6��SS��' $Ӽ��l�J�#��vng�k)��0A��}��1 h����n<EYi7587"<%��Z,�;��R��xJ;K#��W����^*��J���.>��[�����-w��K���>���4�˸n����?$*���/u~{�si���fH�!��0���n۵b-�=�
�<�����L7��^ �ʱb���߱�l	�W�pya��������+�
����`E6jU��.�֐S�R2�2!sƄl����1+ Ta�
�|�C����%����gO�6����v�2	8w�_Ki����/�gSΟL)����IR�s޵��V=<�T��'>����z[3CiBK�' �g�y�o�z��W�
 �ZѤbYf���=�����^�ƽ|��5?|�Wi̜H[�Z+��L�-;�tGTo�����E�u߄wJ�������rI�3Cs��I�LXTY]S��'��Ki��T�%����z,,`�jR�["�*-��GA��L{�`�-�z/�C�T�R��fPv�RR�uG�}k=�ѓ�Px�&�U�[U�U����Y��ki���R[b�K[�R�)�:/u��~��ݾ�P3�ք_���|Yr������?�z�g����4?q[�p!�ť�|K ��}�SH�ۨ8y����l5����5���?���x~���  �IK���eF���!��m/����y��Nz���г�������;�����<�xWP��@��Y󤏧X�+d�RL�XeW��Rk*��tD=^��%��i����������R���f7�Y�t���A�0N��st���6C��P<r�3�X�\� `��X���/�6ʀ���ƞ���P&Fd��N6��],���H��i�������N����������Oķ� ���G��w��~	iaҧ����.˿�d����&�TZ;B<N*�y7��f�M���G�X��+?Yŧƞ]�.�^A�!�⣴�͏Tتe��ײ�ի������z}�Wu����
h"̲`>��Dؗɫ��r�dNإ	S*&/��g�j�(�w8L�qQ.q�p�������S�Ň��ʴ�r�ʧ	��=�_�����WN��i*{-��|���~���r�0��	���	w��^�w�RI8=8�x\p}\���}������Z�ڽ{�ݿ�w�S��,���=,�	��D��,hMH�uB�ɋM�D�o\1e��.�rb�2A�k�+Q����c�i��~�wW�ֻ���-�N��d�x޷$i�95��Ě�sK��wAV��&a�=0�o�{�M�7\!�*)TD�6�(�q�nr�n�r�ׯ<���8����^�_k�
�gk��.tw�6P��2��O��/t~�{��S�[O���3�[���ew@��HE��}�F��7z������~�+XN�X���f`>bz�I��5˼�\�$e��I�i�z�b�E}7P���4�ҔT�����j|k�C�j}�&�,G���ꅔq<U\_/&*����4pݴ��6�c�F}*�����T� �#&��Z�u��Zunqs[|C
ٍK�Q�H�����5�m��
ǽ��vS!T�^�m�ZJ�۾�T.>���.��?�����C�,���#o�R�'�[�@���/�P2�_��SU����j�ai�;[��&kaZ���R����pk5�9Ϗ�$x.�+m?��O���#޾����6�ի�{�+|���k�W���Ҁ�r�um�>�S�������*6PD�]���p�i��~qUP+ �q��;�{�$��}Wn_�zpk��������y7}\���~��_�}��اtwH�����l��t���^���Ջ#ꬸ���)�N`͠�P�x��5�EЈQ�RFk%��u�_b�9����6L��z���X��^~���p��C���ⷿ�{s�U��g>j��`��p�O?�=}j��km~?D_$�}����\?�;�F�|��x�,f8���"g�����Ԅ�i�i^��+�
���r��;>&�%&y\=�]�pm{��u-�+�P�yʜ���M�Ȥ/{�ڏ�o�~��P8%3+��J�B����bG)#s��8�\v���)���xˋ|���?5���Η>�1(	��5�O?��?�aY�����I����iE�I[��XߢV�0�}h�o�ӽ���X#U" �/���i�-��ke�"�
WU������#��W��'�bC)���QR���(�$L����!>�b`�&ȑӄ[��ؕ���jŔn#c�D	�/���~�ٯ=y��������n�����ҧ_���$4��sϾѷ4��B?�a���{
����an3Z[px�����{���%Ǉ/��J��K��Z�k���bAkC&��^�M	�
�B8͋�N'@��i3/W�Zsx�����F%\�I���+���'�9#%B���d����)���pLލB��Z�l#Y}��	 2��4ٰ�4������k9��J�WA����>���8��-��7�������@�/|�ؽ�i\��h�G�y�����^�N��wf�ߩ�h�����Ui{�Z �Td��^��G��7mܫ��#��f���a�
}������J׆������,*�#� jC|��I��WhRQ�u�K���%d6�f���i���U����\���w��;O�}�c��̻>��/}�ݓ�s����p���7�6A ��_�E �VA�3�y��镯���t�.>Ȍ�6ײ���{ҖI*�r�2� ���s�>m�P���ٔ7��@��xS����]�>�
U�b5�UKIu�����e�i�GǞ�2��qA�x��y+RE`���{ΩW��(/�r?O��r��/Q��H��r��;���/E����=�;��O���`y������SO�vz[m�gAx*ߣ��Է�ջ"� �C2IUXUX��h��d5�㒮��R���Ůq4%+a����{�}�EM`B\���� �����MLPb7MP.>�E-4�4�\�����������������O��,������e���[Z��?��O �^�����>�j~��[o� <xG=]�u��
�>��{���і;m^��T8^�Z5u����54��mmV5�&�'o
�v�k�z#�����3!�U���(q#2��ܵ!o(��p�˔�g��I�.�,̩��2_'N��k����?���?���^�� ��}��F���t~��[��?�ҳ��P��׸x�S}����[h�Ro�N"����P}Z���[*8a�������խ����c_q��
���7�.?IB�,�m��*����>�0��וf�����m���5-˂��Jɨb�1S.Z�W%O��������px�s���/�{�ٷ�-�<�����o�� �g�ԧ���x�|��� rxn�,�����6�<S8�J�U��o"z��o�N�Ts���(��yO
�jz6O���"������
�6C����ܭ-nk�$))aۤ>�i�2"��2%%NB����J�f%>�
����K�ӗ�����qY꧙���F�^|I_��R�L�Uo{���ѷﷄfw�/|�v�j5��@� /����#K]�&�h�Y[M�IRQ6�g"�邈n�-�iOL;UL
ͤH`Ndc���X��J�d�G�*T�`�FB��5���B}�+��De�8-3��#�*�2�~�'�V�J�����<����������O������/�u�4��|��ѷ"�JT�}�8�M����p��~�N��p:ͻZka���:�D�ۙ���������nI�Q�h�k�y^��T91133)"�b��f��@�Y�Z�\r΀���W��X))1	@ں�-�1QQc�
�
�3���9�gN���U��N���,���>+���S�S^��N������¯��'�
�����w?�Y�؏��}�� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��1�Ӓ������   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X    IEND�B`�PK
      RZd��   �   /   images/a262aa33-74c4-460b-b0ad-c746896f6744.png�PNG

   IHDR   d   d   p�T   gAMA  ���a   	pHYs     ��   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X  �IDATx��{y���u׹���Z�j��ez�����L�b'������2�eH$BaJ�@�dC��`�@��![G6NlϒqO{2��=��RU]{��ۿ�����1�'��n�u�{�[�=�s~�w��ʥ��1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�l�c@�a�z��Ti�R��)�|�H)����]ǧ0�Vg�¸K�F�Z���=:0��y��8L^a�&����4�"ϨH32ʐv4������>Y��6����=�n� ��w�H��)�~�����t�g��!�<T~V�Yz`�����j����ר�����Z�:@N�NF�ޢ���,S�ޠ��NY<�Zk��J��� m
& ̡T�nW���]����{}*f��>s���m�ݽ㯐[����u��)h~�����>�����R����h_�М�NݴC͠���ޘ�g>�?���g�~��P�R8葉ڤ+�T�O�8�,�`�UZ�	!�n�6�a���y6O"ǭVk��D o�D9~G��[�m���^�u�'^"�[^���O�N����+ DF�u
��v�����/M2�P���&���8\��
\��w�z��V�K3�K3���h㇟|������~ݟ����W���f�ȉCD�M"�!Y֕�.���n�Sf�	ch��G�&�q�H5���*o/��%�ݼIj��KI�Z����.J[�(�\ׇGk2�j�4���X:
A�tԿ�M?�Yg����K_����pkC通K�23�*0o�g3�$����0�v�g~�/+�W7��|��ּ�,un_����� I;���\��u��_},�~�n@"��-ob+b�v��X�I��f�L]�Һ^��U�8�E'?vV�x�C�k�;���M�}$�DLi�S����mQ�Ņ�:��(_Ug�����F�����	��ġ`VcrDqf*��q
4SU�NLm&U^�������G��i�8�3�.�۩.tؙ9|fp�[�D����W)�lSg}�����ѡ��0���%�]���pa�[���>PD���~󧢵�� �v���ԡ�����?�j�UZ��ε��@��_
��e���,�=McB�'�pt�&���.���
{^�K�zst���t��I��#���\N������r���4a�8&:��i�M����fS޻�0�*N�� ��%
V^��'B�%���w�1�@��Yuh$L�wQ&�0�3��	B8f��e�wA���Hi��%�?�p-,$|M^�0$ln���ÃN��'���S���;u���}���~g�| ��eP�>Gӧ>�����)3���I�+Q$d���򼴍�*ձ�aѣ�x�M�"D�ܤ,=E��Cdẝ��HKb�=~���kur��0!�-�)���!��D��)�px0D!�`����!��YҞ+sU9��x�T�J�,�OR@do6v�"�J��:������gB�K���E�����Ԡ?±��� ����s�Kh���+��7^mn����&]
wV�:{���i��u�Z�|�I��'��&��=�{��֠}m�r�<�r � ��c%ED��*�	���8k�0�Z��5�׃S�w����i@�g�ׅ�âz��w[�D'��I�Ar<��a�L*�އ\M����G�+�+��߰s[�����
��T�l1�z��=��.� �v+r�v��[�D�KO��c�	�K�N����[_|���S\�m#$ł��y��s��~)�oR�"�qm�ߵU�/�ԃpw��
"��U��2��Nڦ�<���w]B�^�X�U�F�ozZ�3d��(w�m����&�ҳɂ�d^J��)$��D� ]��X0�*\KIy,`Z�S�oا\G�څ��k�ԫ����G(4ED�+�i8���\r;Y_�Fa�bn���V�`���܉'�n��z �}G����#7��{�B���/ga�`:��v!{�%Z�A�q�P�w���~CYT�UM@u�C�D&�����m�O���KY`��Cs5�e@Q�f�\Z�m��-�%*$4�H`ٟ�i2WD�L]VCq�)�~�dQE�:�)IX˵喝
��O=E>U�)��:[[��Bβ�saȜF3�`H)E1��>>CN�?оs������=��;k�.�$�ҩ��x�~���p��_Α7�p�&q�@NTNu����	yф���ά�K���	]�WQ�6���p^S7����N�z��7e�WY��G�95�F��+�ÁBሚ�t�D�,UX�/��p $o�T(M{5�ր�2�gBrNa��r����
�7_׃s̟z���S��\!3X#߳�7��0��p�3��<��D4��Y���b4~�:��˝�7^�H,P��J�ܰ�K핛tv�y��'�w���y�����a2UNQ��8���/#z��!X�4Ee�w�.���9��� �ޙш���.U�5rI?��H�>��!���~�
S%6Y!
F��[ͪJ�亢�"PNтĚ�Ҿ��\�*Ȫ"�윬c�*#��%j��}���y�����﵌r+���Q����5��#w�<� o`Nٰ]M�꿞=��3������i#$�z,�Sm��}ݕ��}�{���ޑ(P���̄ZP^U<P��7�E�)s��p� �Jg�"L��s���8=�8�&Q&	�A@����d��U��Z%p@ e�w�C�� jT���xbn�[惟^��.�ӶxmhI�R�8��X[;��Dn�E~�^��WR# j.�5�RX�_�r�+��]�ʜ-��"���^�t늬դ^��G� x�s�⿸���ԉ?��Q���:�o��� j���g㝫���8��/�(���E�a���r��j�Tܻa/k8S�PY$����I:9s��;��1�M��0RE��<�Rھ��DR�y�2���D�*��$�ETdF�(�8*4�uD)1{6G�����@]-��=F���r��q����0��؜(y�s����@onm/;1�y�&�'����YH��.�KT]xP���SY2�A9qE���	r��������������έ����{>�����@S��/�c��eu��ʘ���	9%�Qڪ��x�"�4a�$ۡN�o��t���"��Z�m�O�ȉ�/SmΞ���%���b[�Ap�����29?gi�IH+�� p"��� xH_�\U�#�8 �=���� �Ʈ��Π�P|9�G�ex����)ݥT�$��5����)L��H��=�c-9Q��3�C���"��BS��4�=w9Z~j;�~����i�ě�}Ű"a��$�ڝ{<��X�1x;"g U.�*Y-���$�0��=��FG*��wi�f���zK�l^���~M��!t`����E�ޗ��5@���R�3�7(T�rl��<��T��;D5�PD��ѹ���d����\�p�!ё�I�#&��Hn=�Afa������[�M�����ox(�}��jߑ5*8�ҷ��D]�kduƵX���E��e��g���s5��w: +�KaS��q��0Y*rc�dZR��+J�*�G�Zc���"4A30��7���ޯ�Q�/�޸D���xs��D�p���.a����6�9%�3ա��XYn�"L[�˭"� �� 1��MR��(a�F��Pcs�6���w�UD#�ƴ�k�:&g�ɻ��P����]^[U��գ�W�s�%���@X���f�S�?��:	���.�B�r8�魐��57�ڛ'�G�͢�k�$�\.�Ӳ3�������|�R�|�|�܁�ڴ���P-���ץ�+Qhlo�)�^��˹!;�S��1C'�aT����Uz+�t�$½�;j�9�d(t��x����m�0H�Հ�"�Yi��BT������5���8R��/6�̽L�FKn�M_r;4��<�\�؊K�E~�%ut���ص;�2��e�@4�����*kY4S���X/���9������
�Y
p=���8�8,Xp��ͽʶ,�{F�>Q�H�Q�Ĩ�SCsnF���g���T���胁őX���}d�$PJR�_Ξ)�
���֠�hGh[���j����'M1��'�>�Hd�D5��8R��,
k"�Y!���C��\Ŕ�AqY�(7��=�b�H�Kr6���e�Nو+_2Kc�����]9ڪ�£���a�Y)@+[3N���?�u@Y�I��2�a^I
��a�|&R��e/Ki�Y����������<}8���$i��{{*2m��"��ZjF�R9\ c�YZ���V�#�j)y�*j�Pj�T))6�����Q�Ƥq��(؟���Z�K�כ�ό��bЃ�l%"w6�s9j�k^\	�m��J� ą�|�(�MҜ[_$9��.e�h5e��ؾ�eJ�F�M0>ߵ�����C���W��4n�&8A�{�^�U,|^x[]��~{�/ۓ��S���r�*��VM:�Ibh*,J2�{`PY��-s�&BU�S��!b%f6zx�"(���u��_NM��ϯ�]	p���[ِ�������C(A��ʚ�&V�%n��Ҳ��m��XZ)�77�lH>�~X���w>�ⴇ�P8Y��e�z��>�!,�S�}%�[��˕�P$+!g�0��Qd�F��-¬��X5�@�iPE�vٟa�T�r7����hޅme���-�a�����Ɣ��;GМ��`��?��{��~�ɿ��'�������C�r.r��Hf@�޾�ѹ���J�ƲЛ�J8����1��� B.N0���=6ۈ3ei��0����E+<÷�V�sI���ϋ{=)�[Q�����#�Ap$�r��q�a(�`�FQО�Y��jî1��X�~�ʍ����C��V!��e���z�3�r�[)W�`�'��?�%��_x���gg�~�Gk�7l>�UH��E�ǡ.J!�dv��:�Ք&�6N���&�1�Ri3צ��=#*�!>�
�mI��P�{�0$j����쵲�ABf�Y֒#����j�����K+GDA�iy_dv�Q��M��T�b���xm.��P�vű|����g�e�X:�JP�W�})B����qQ���H��=���t{��?;�U2�1�	���`���'�~?l.���!Q�w+gD��w��<F��8� ��#$�I�G^�Aa)�un��-O!
c�	����ԋ
�	i(6;��R��	�����|#M�RJd�sRa��
VO^'ANL��Y�k���PY��6��Z��<mMf7�4�t&{,E)�*v�t$F[��1!,�Y�y�s������}2;7YW�����c�q�u�x��T_,.y�}?}�y��,�Ӱc���Z��团�`����)&��|,Q�%�3�Z�T���OD�R����M�όy����|DJ�s�<���O(]��Yx�L�|��X�ǀ�ANY�ؘ 2��H0/n]��z�̍�s�B$+D���"Ys3�T�
Z9?�`NY�h$�(ͲQj�cIQe�_�)��T�~.�t�̳�z�U:�����!�����(��+/�����_s���n�E}��P�{o�����\P���r���J*@S)GG����Ae!ȋ�G\^���P4l�ݞO��+�;�,�}!<��F�R�L���=T`��v������[C�����8/QV�I��@�[�%���-s"� d����uH2��<�P1��:h��gI>�b��I�ѯ�Ch5�������7���st�]��\�v�~7-_x�K��c����YtH��O�-��:�F�"iK�\Ŀ�׏���4�ϐ�x��
�d���Y���Oi+���V���!���h�w�e
 Ң)�;�YِR;@nom��@O���#&���V��UBq���ͯE�.E��4�΂+�5YO�{�F��`d�mp_>��A�Q/���t���h�(��;�_�Ï�|���|����k����W�n�u�1��H꿡������H1��;�^�[��dQ!G��Ȇ2�@qN��A!)�k�ҶVE�V��u2��f�u�k$xn��(0p��]6�F�DSFF!^���+
��l��?W�yn��\Ԡ)v(�6�r�u$��k�
PEO!���$c��'�,]
�Q=�st�t�\���ׇ^�������yo����G����!�v@fg��k/����?���������S�ҡbЅ��e�~i+e%BVG��b�f�n��Cb,�N�w���Ƚ �T�k\�K��'���V��h���]�B�� ^�>]�����lM+�wJ�2u������5)Ly�2�MR�UI5�}��L��k1����k�	oN9Vy�߇�#Y1a;T�&�.����í�~��c������c��i���?0��e|�)�u�T���[itď��FC��'�Oūx��i�\�s����3Μ�-���'���*��jו�6$���-��4��"k����z��J�Z��sը�Pvo]B5��\Q�{߳5�[%g��ٽ)8�eC��0�,~F�_�J��@t�4U�*(�R��#��>�M-�hQ�3�܀�t�m�e�l�a=^s��������~�wx�̇�w�������K��|�vV.��}�?���?b��;����"�e��=�f/.��kT_���En��u:��!j֏H����V��|W;^�K���MD���*��4���AUy���Ss)�f������|��#;���.�u ɎHw���.!��#К��BZG�����8�%��N5O�zGSY�u'�}����O\B� ��Ȯ�H�N���a�'.j�.Ҝ�g)�#p+Ti-Qe��E����a{c��n.�������ճF��w6�S'�������:���H�}R�sn)���>���z�&�3�Uϣ�?M3�����Go�V�3����W_s+��&��N/�G�+���Q���Yz���k۝f�f�����@{��㙄�"����Ju��9�r�i�v������������X��� �:��LT��N{�/)<L����l߭;�f�y�5����ߗ{�<r����.��y/��^"�@�ZI=�F?s �<8^0��U�s���t�s;���H�}oJ��y�V_y�q�����d�����~�v>��n�%G GS+]A1��4��x*�������D�ۊW�=W��k�>��/]�򯷛G���	��P�_'�*�.kqgv{��RoQ7�d�*qR
}EQ��0�і���|�>9Bൕ�e2�-�i��,�bؕ=>'K�w6h8�KG��� `<PRvP<�)���y���?�ɠw��G%�:��=SSt�0Eu�婙�H�Z��S�z��M�yם��?[�N����s�<E5�X�����w3���}ȁG�CwΝ�J����is��*4������V��6}���ȼ���T+�����ڌ)	w�9�_����W~��W.�C��%ZlP-h������}/^�L?N/|�b`|P��֚l�nܜ��U�y�ؗ��ڇ2�[��}�[����<t9`@K���w:�W_���BՇ�{典H�o�4�f��2-��_���[�p�C��
��9.'u!\1���tz�5|�|��>t���W�9��D<����Auߙ'�~�s�"�?�7i��D�����G~��_{)�]D�D��.
ɵΦ��j[Mz��ץg�͆t����q����r�N<�m�W.~���CTi�݋�%�W�ƉluKu�P����FS��5����� ~i�~��wt�?�}�w�����O��O���wf��c�W�c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2f�D�{��w��    IEND�B`�PK
      RZ+L$��� �� /   images/d8ab57a1-5a79-4c55-bee7-02b60939cb6a.png�PNG

   IHDR  �  %   ���   sBIT|d�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<    IDATx���   �����
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �ك     ��FPUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU&��M    IDATUUUUUUUUUUUUUUUUUUUUUUUUUUUa��c-�
�����>�;o����y�G0�Nj��I�$ĎZE��J5A�04�q�#16Qqm5��4E	j�T
!!����f ? fl�}��>{��?R^*�c33�>>���Ց���?�^?-                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ��,�     mߔ���|>�lGh�ݡiFuQ��e�]�!�˸=dM^�0�R�41�bS��&tR��,Ƽj� ���:��w��i�BY��&t��Y]�~
����b��jR�T|�"�e�)}����<̿�{��i��9k��f��,�iBj�,Κ���<��2e�<Ka�Ĵ,b��&��NZ���N|8��IȲIȲ��Ms�A��x|�T|?      6w    6��M�E���ٞ<�v.��3��κN��&���V�:����R��	�:�~J�h�ԫ��KM(�&u��q��Y\�,Ty16e�e�<�y,�4�iR�汙4Y�Vdi5���ңyjm�x<f�ñ��4�v���     ��g�   @k������U鬦ΞR�tFHiO�⮐Ҏ���U��7)[IM�u4M,��?t�9[QLE�YfE�1K�,6kyOĘ1>��t<�x��CY�|wQ�#������ش]     ���   ��暃)?������9���YM�Λ|�2�ݩ�;�*�Sؖ���\�aUǁ�:�WLE�f�"Lcֲ�Y-��x��#����Xք�t�pd�ɾ�г{����X�]     �U8<   �q���it���9u�zz��c�ϮR<3�iǲI��*�j�l�r�7)em��ɔ�aQ�a���G�<ϲ��e�h�GR�{5�g<�G�n     ���   ��k���//.
E���鼦i��pf��g,봧��e�5u��
�]��eQ��<O��<+������,�V7���<�{���߸     ��   lb�����a/]�pQ��y�
��M<�j��zvUu�qN�,��(�4��Eɳ�P,·��y�����߿~p_۝      m1p   ���㵳VcxNȊK��paӤ�.���*�S�*�]5��v#���,��"����X���y^��쾬�ݓ��e�k�q,��     8�   ֱw�;�<\^\�pY�l�Q���eϮ��Բ��h�T���^YM�W�y:���N����o���k{�1ǣm7     <Y�    -{󍫗-���y���������:���6�"�N'>�)�w;��@ҷB�����7_׿��>     ����;   �i0����sBV\�\��*\�(ӹU���m��b�nN��H�h���쾬�ݓ��~����      �   N�������/Z���Ԅg,���e�*�aO]'7��Z��y���y:���}Y7�������싳��     ����   �	��SW����,�p�r�\�,���˰;%�[��%���t�j7OǊN:\ᮬ��S��3��ྶ�     ��Ł+   �c��ӧ������uxfU�s�2<��°�6���ۉk�N|0��;!���Ν!�6�i�     ؘ�  �-�7oN�8��04ٕ岾tQe�W��E�v����yXt;�h��-�pW͝��?=�n�     X��  �-��[S��gW,���MJ�.��E�^����4ޓ �R1u���n���)�����~�|�����7�e�u     ����   ؔ�z���2{A���ez޼�evvݤ��6 ~ �b�)�#�n�f�I_�v�;�����>�v     p��   �u�X<w��\����/.�pnY�neؘb��N�����N�Y��hT}����j�     8��   �[��?sѩ~�n��e�t1�O��0l��S�ȳE�S�wý�n�rȚ۶W����ش�     ��   ��������U�mw�~�����K�yﵱn�     x��  �u��7�^�,�W5ux�L��e~NU7��� �x�<.��x�Xޝ����<������j�     x|�   �i7�)�q|m��Jً�e|̞֬Y�͎�� ؼ:�0�v��n7~=Ϫ/n˳��p�����     �e�   �R���mۮ���˲~nY��Uܕ��{	 ZS��v�ov���a'��s^T�囮����     `+s�   �T����ű�^V7��yx��"\����� �'��v��A?|�׍_��������     [��;   �ǩ�Z̮��xUYƟ����E��� 'K�&�^so��T�����_ܲ/���    ����   �{����k���*^Y���f����IE�] p�dy\�{�^���ݩ���8m�     6w   �1����wBx�b�^:����evf�� �!�n|�׫{�������һ��&     بH   ߷����:��颹b��.]�aO�M ��t:a��5�v:�K�����4��x���     `#0p  �-��[S��G&/[��˫e���<^Pա�v l6E��A�F��Љ��x�ʧ�{m���    ����   ��k����f/��xլLW�g�%U���4+�Xz�p�n���G?k�	�w     �[�   �I���`�     ?`�   �Ⱦӽ�e|�r��-�Euzm7 OL���^��wXd��v���뇷��     ���;   l`o�/���y�yv�b��� �\E��~sϠo۶#{����}��&     8U�  `y덫{����z�t�=^Ƴ�n N�^7>��Շ���S������ʑ��     �d1p  �ul��#�z׮W/����Yz����!y� B!�Ҡ���4_*���l���n�gmw    ���@   ֙�7,��\6??+ӕ�YvYU�n�M �Ɛg���}�^���W��wV>�v     <�   в��;�W�����<aY6;�n 6�^7>��Շ���S������Ѷ�     ��b�   ��5S~���?����Y�b�Ȟ֤��� lnYM�5��u��Ç�5��{��u�]     ���  �4���������gg����e�� lm�"�z���~���M���    �z`�   ���ϛ��5�<��Mni ֥C�u҃�Q�L/�>�=�>>Ǧ�.     �w   8I~�wӎ�._YΚ������2lk�	 ���a�?h���O����ۯ�~��&     �w   �	���]�6˯����<]�4)o�	 �dʲX��"~r��{��o�w��    ��e�   Oоӽ�e�+�Iz���LM�� �2z�pl4�?���C�����ql�n    `�p    ���N�o._]Κ�'�슲J+m7 �E��A8��U�X;x�MgM�n    `c3p  ����6�0_f���t�l�Y7�h�	 `=+�X��A�� k���h�	    ����   ����t�٫'�^����<^ؤ��� ��R�����_�Y��w��_l�	    ����  �-m߁��e���t������MM�Y �$�uñ�(|��U��wV>�v     �C{   ��k����N�Z4�?�N��,ʰ��& ���׍�����y߮0��x���     X?�  �����=�L^���-���0j�	 �z�pb8H�Y���~��oxC\��    @��  ؔn�5u}g����~��4���°�&  [���h����=�ţ����h�	    ����  �M�GF����6j ؈��    �.w   64�v �ͭ��|4H��     [��;   ���Y�}���k���Mf��u�zm7 p�u�8�/���}\:x�{��u�M     �\�   l�L�9���vS;  !���ĵѠ�\Q4����c�v     ?9w   ֵ}�{�Ez�ڴ��r�V�� `��v�GW�۲a�Ͽ����m�     ���  ���;0ݻXf�2����e��v  G�����B'���׿��     �w   օ�7,��(ӿ�L��拴��  6�CZ�o�{͟w����4�v��&     ��;   ����Z͊1��W�-��R�xN ऋY�����m��Ѧ���;ǻi�	    ��p   ��j��#�r�ʵ�E���i���Iy�M  lE�-F��N����4���8�m7    ��   �r�L�9������NL�U�m7 @���p�|��I�}W~p<�M�M     [��;   �̾ӽ�"{��$�tY���{  �t���h>ى�}��Ŷ{     �*w   N��x��!��4�j6���  OT���F�/vv��p����{     �w   ~b�ޚ:_{���ɤ���4NӤ��&  �I�,ԣa�~�y��4���8�m7    lv�   <i�L������I��U�m�  ����ĵѠ�\�����m�h�    `�2p  �	����.LU�׳Yx�|��v  �n�~z`��>�+_���x�H�=     ���;   �뚃)?���5�I��ӵ�MY�M  ж��z4��2��c����86m7    lt�   <�7߸zY9���Z���
��� ���[���Q�W۷��-�;��    ب�  ���5;v�v�~ym�]��Ƴ#  ��Ŵm��1Z	�F�?�e_��]    ��)   Ba߁��r�^����ê��{  `�����G������'��    ��  ���޸�g:��Ģ�'�y<��  ج�px4h��y��[^'m�     �W�   [п=0}�t��գk�Uuzm�  �VQ��b8�n������i�    `�1p  �"��?2jv�|�d-��Y���  ���txǶ��^���7]m�     ��   ��o��T�򍫓�eU�m�   ?�Ӊ�m���۷��-�;��    h��;  �&t����{w�������Y~ij�  ��Ŵ���w�Qv������[��]��0`V�/	[X��-��3͸����,d#l˺�lac!�<:	�f&�C҇3a��e�t�	`��]�/w}�g�H;!�m$KUO-���R}���.���z���P���N�����g��E     K��  `�hW�١Ο�����Ƒ�=  �S�ds����C_������    X*�   +�#������-̗_\�XJ�  ��R��w����n�k�FV�n    XL�   +T�O?[�ϗ~�Ӊc�{  ���_C��^�ߴ�����{     ��;  �
�e��9����˯.�XI�  ,��������3{w��<u    ��d�  �lnL��b࢙VxG�OK�  ,�l�@=���s3�ٳg�|�    ��e�  ��]����.��	o�塖�  X�*�02���j����W��N�    �D�  ,C[vΝ�lW.���^^�XJ�  ��R��w�V�߽�1�S�     �(w  �e��?����]�����{����=  ��V�ŇF��/����o4�N�    ��a�  �������X�ha.{g��S�   �K5����P��m4���    x<�   �\���W��f�JoȋXI�  �n�R����H=��ɫ�K�    �Gc�  ����X~�=�w�����,?/��2  `�eqp��kh���n�k�FV�.    x�!  �h��'gZ�=3����	R�   �B��?)���56̤�    0p  XD�]�:k�.�h�F    IDAT������c-u  �������P������^Q�;u    �v�  ,�-;��i�+��g//b,��  8�R��w�V�߽�1�S�     k��;  �)r����C������d�R�   ���z�70��>����Ȋ�=    ��`�  p�.���\��əp^�֧�  8�j�xtl(��H�{��uR�     ���;  ����3f�}��gK���š�=   ��Z-M�_���ܰ-�N�    �N�   '�#�6��ٖ���<��{   �R��5���F���w_:x0u    ���  ��׵_�l[��Jo(�XI�  �R��uG����t���#?J�    ��   ?��]ͳ�م3��1��  �I�R���>X+>��ꁿI�    �l�   ����;ڥߙ�Ϟ��  `����`q�h��mώ�o��    V&w  �����8�����5[��{   V�z->48�a}��F#+R�     +��;  @�ҽ��͵/��	�;a}�  �ՠ���g�a�追��:�{    ����  X�>�{f�L�o��l��;�8��  `5�VKӃ��ׇ�=7l˦S�     ˗�;  �&}���ӳvv��\��^��{   ւJ%,��?�0�}ckv,u    ���  k�%�7��5���΄��  �Q)e�������<���Ȏ��    �w  `M�����|q��l圼���=   ���=�h4���    �3p  V��\�|z�.�0l  X��   �G�  ��#�����9�a;  �����}d}h�t�`�    `��  �ʅ����b�a;  ��U.e���޷�   `�1p  V���y~k�o��\���   �C��uG�������۷����    ��;  ��]uS����Ǧ�7�"�S�   p��   ��a�  �H��   k�#C���]�F�ǩ{    �S��  XQ>�g��3S�˧�Jo�E4l  X�J�;:h�    ���;  �"�  �/=2t/�g�n�^�/u    p�� �e�g����ט�-������  ��TκcC��#����K��    �8w  `Y��څ�L���S��s�"VR�   ���KYwt��퍣W6�f�R�     '��  XV{�������ү��?u   +O_%k��o�������f6��    8~�  ��p��X/fZ�N�d��za u   +__��_^j{����    ��� ����X~�]�OL���t�h�   V��j_7>7����hdE�    ��  I4�4Sn�?9�}�݉�S�   ���kف��p�MW�%u    ��� �%w�u�s�'�-�N�)u   kO�(>usc��S�     ���;  �d>v]���3��f���-   0\����]77��"u    �� �E��څ��-�mss���n  �.�CC�����77����    �:w  `�||��''�W�Ε^��   ��R��p�Y_��4j?N�    k��	  p�]r}��|��rr��K����=   p�J�;6�������F#;��    �w  ��i4��������윢���=   �DUʡ5<�����u�of�{    `�0p  Nڭ���/��NNg���0��   N�j%̍��/xa톯���{    `�3p  Nʥ׵ϝ���7[ac�   X,�Z<86\�����    V3w  �	ٲsfe��BxF�   X*���G�����C�I�    ���;  pB��n=wa�h�̖_BtO  ��S
�.��8�v˶���{    `51F  �����X7�wNOg�SQ�J�   H�R�Z�����S;���4��    Vw  �q��+����/��>�����=   ��T�ar�h��F��;��H�    +��;  �.��}��T����NO�   ��@-��v��Q�f�    X�� ���k^35��[Ȟ��   V��T����)��a���R�    �Jc�  ��ˮj�5���s����~   ��R)���|������ٱ�=    �R�   �c��х���ӳ᝽<TS�   �j�WɚC���N�j�����    �;w  X���X~�]�OL�:�0��   V��j_7>�w{�3�[    `93p �5ꣻ��99[�x��=)u   ���p��`�}����    �#w  Xc.��u�\>1�PzE,
�   ��JYV���^�]��1|$u    ,'�,  �F��������u��t�7zE���  ����/�.���k7|��,O�    ˁ�;  �7Ν�+}��	R�    �\�nͮ���ڟ�n   ��� `�ܘ���N隹��KS�    �'��C��#q�-����   �T� `��1>R��]S��Wbʩ{   ��S.���H��KϨ]s��Y7u    ,5w  Xe.�9������N�M�   <1�Z<<<P\wKc��[    `)� �*����.�_��J�   ���T�����.��#?J�    K��  V�͍ɱn��~�(b9u   pj��Ywt$�i}~�={6ͧ�   ��d�  +T�K3���cSჽ^H�   ,�j5L�ǽ��1u    ,w  X���l�3��5����-   ���?Z?�_vö��n   �S��  V�+n���x�S�ٛbt=   kU���FG�7K����fR�    ��b  +�wľ;�w�������П�   X�}azt$�zˎ��S�    ��`�  ������s��u����-   ��48�qCo�'�� u    �w  X�>v}��_���L��E���=   ��V.e�������\���r�N�    O��;  ,C[�i�ob*��酑�-   ��R��o-7\Y���-    p�� `���YsE���\xe�   `%���p�7���/nl͎��   ��e�  ��{��g�������}�<TS�    �C__��0>������-    p<�  ����gOΆ��VvF�   `u�wm�ػ�[���    ��;  $��19�˫7LΔ��ks   `q�KYod4~�:ڿ�-Y3u    <#  H��s黴Ӎ#�[   ������6����ڟ�n   ���  ��eW�Κ�������-   �Z�ő��o6��_�ؚK]    �0p �%�h�����>;]��^��{    B��/�o��{umo�    ��  ��]��8;[��يg�n   x4C�J�}Y��S�    ��� �"�ژ=�٫|rj6{S���  ��\�z#�����m7mɚ�{    X��l  `l�����Bis��R�    ��z�tx�@���F�[�[    X{� �j4�6���̖^��   ��*eY1:\���Jk�͍uS�{    X;� �ٲ�u�����^/�S�    �
�j656��y{����   ����  N҅���쵲[gf�KR�    �jY��{�iC��Ɩl"u    ���;  ��-�Z�Ofw��   �rվ0=4R\{�����n   `�2p �'�]�gw⭳�ًR�    ,�GNs_7ػ�W����   `�1p ��eW�c�%�<�R�    �P�����'n�f�˩[    X]� �8}|��Ǐ��:��I�   ���xZ<���S�    �:� �O�h��dhm��*��W�j�   �夯/̏�Ľ��>u    +��;  <��]?�����-���Y�[    ����⻧���j`�    V.w  x���>1Uz^ľ�=    +A��F­�6j�M�   ��d�  ������̵*7/,�g�n   X������G�o�V0u    +��;  ��F����3ӥ����   `%�����u�s{���M�   ��a�  !�-�.�nz���يg�n   XMF���*�x�����R�    ��� ��5�4Z�&�J���v   ��Q�d�u늽�l��^�    �7w  ֬�nj��С�w��3S�    �CC�wϨn4��n   `y2p `Mڲ�u�щ�9�C�   ���Z	3�C��[��?S�    ��� ��4��C��gg���S�    �UY�ǆ򿬷�?�gϦ��=    ,�  ��^�|��t�N7�n ���O��NߐUƧbob*�s��E�* ��z-�^~���o�n   `y0p `ջ�1>R�n��+�)�k`  Xd�o�_xm�?,���gc>1��"�����lȍ�!�R������ѿ���n�    �2� `U��1��cs}�۝�>u  ��r����h�=�3�^7ƙ�����c�7;L�ְz-><<P���F�;�[    H�� �U�шգ�}��TxG��{ `����C�e��7�v(�fb>1�ɩ��O�^��b5��Tʡ�n4��-����-    �a� �������N̖oj���-  �V��E����N��i�B~l"��&���ə�G��z�����@����R�    ��� X5�X��mS��ʋxB'E  ��S6e�7��<t��߼qz&�G'B��D����N;8�`���º���[v�?��   ��c� ��p�M�:T��B3{f�   ��J�����HX���qn.G�b��x�ON�|j:��3XB�C῎u���#�[    X|�  �x[v�.8:6�y�O�  �����<<:�����ڡ���S����d�&� +Z�Z��0������   ��e� ���h��u:����/O�  �k�|Y���3����E���wt�ȏ������1u ',��F�����]pӖ���   ��a� ��t�5��NL���v�`�  ��=��Y�k~������L���CG���q�w���V��6��͟�j�oS�    p�� ��4�z4�o����Bt=  �X�J�xse$u�OS!�?r��x���"O]��)����h��O�oO�   ��e ��qō�>Z|��ʞ��  8>�xse�^��'"/B���C�b��Ѣ71�X������Q�?�hJ�   ��a� ��p�5�ߞ��.��؟�  8~�}yy�̧d��'#�C��2xX��}�̺�x�M;j�H�   ��3p `Y��1>R�n����N�  ���<#���%���R����w�h�;x8���`��X)ˊѱ��#/����s�<u    O��;  �֖��s&gK7�;q}�  ���Jo;�<��c15[!�(��.�G�C/�c�$�5k�����>|㵵{R�    ��� ��4�t4�vNM���XN�  <qY)�w��2R��RꖥP!�O�ށ#y�ჱ;7�tw��V�dͱ���[w�� u    '�� �e���S[��s����S�   ����\y�ɧg}�;Rh�B~�X�>Z���n/8�`	d�R�����v�M[�f�    ���;  ���]���d���š�-  �����d�/{A���#�C<6z���'c��	`��U㡑Ӌ߹������   ��c� @r�F������;bt�
  ����Y��ח�Sw,7�X:���Gb/ϝ��*��36�������-    �t�C  $u�M�:Xܱ���L�  ,��»�^-�<�~,E��d�8��x8v��P�nXm����T��iI�   �c�2 �d.�����D�5�C�  `q���*��m}�;V�,qr:����bw|2橛 V�j�4��uŶ���Y�    ��;  K���H��ur&;;u  �4^�R��)�Rw�D�V���������c���pRJ!���7����W��|D   ��� ���^��ډ���V+;-u  �t6��U��s��+]��CGb����{�P�u{!�nX����R=|�3�ڏS�    �O� X2��no?:��PN�  ,�J%d�z[e$�<�>Ub��D�8��x8v���lw�T���F���j�    ��	  ,���#������d?��  H�o����J��(�B���C��bwa���xeY�cc��G^Կ��fy�   ���� �E���:2Y��V+���  H��/.��zf�?u�Z07�����ٹh�p����6�n���S�    �e�  ,�Kv5?49Q���   <팬�u�(��Xk���__�=}}���+k��   `�2p ��ۺ��`�6��ə���-  �����_ke$FϦS���{љ��� �"+e��h�O�oO�   �y�  �)���3ϟ����B+{J�  `���_��r���~����m�X�`cK6��   `-1p ���|m��N��+{y��n  ����l����f��;��fB��y�����`����j��8R\t����   `�0p ��qG��������!Dט  �cz�Y��/+����eY��1p�ܿ?��!�nH�\ʺ���n�5pk�   ���� ��r���3[��f��9�[  ��ox(�~�*#�;8.��x��{8�>t v{=cw`m.��������d��-    ���;  O�%��wL�Vvw�q(u  �r��[*#��PJ����uc<p$t:Xt���X�.H�V��Nۘ�mC�K�   �Z� p��X:[;�'���F)  ��yë�OٔUSw�Ĵڡx�`��{��LL�<u�R��Ckl,^w��S�    �F�  ��ƞ���x���·��n  V��>+�����;8yss!߷?v�=�w���\w`��J��n����<u����Ϻ�{    Vw  ���]ͳ�Mg7w:a,u  �r��7��2���S'�B��������n�b�&��00�鉶��L����-    ���;  �e�5�-G'��ɋXI�  �lY)�w��<Z��<�^��"��b�����������r�J6�n4~���o�n   X�<  �q���qp�ݝߛ���K�  �g��<��Ӳ��,�V;쏝�(:�s����Uʲb�h�چR��F#��   �$� �>v��K�MT?�lOJ�  �./~^��E���;X:S3�w߃yg߃���!��XCC�w��X_cK6��   `�2p �Q}t��;�N�w��0��  X}N�*����P��^��C�C��}Egb*�{ N�Z-]?Z���+����   `%2p �_��Ѽb|"�`B)u  �:��Yx��ˣY�9�Z67�}�c��N��Tw`������pw�m�}9u   �J��  �h��C���c�~z6�:u  �������cY%u���ñ{�E��؋E�"���e!�_����[    Vw  B!l��z��T��f+;#u  �6�̋ʵ�=+���`y�o����E�����B0uV�����GG~�m�t�   ���� �p��֯N�d�w�q0u  �v<��Y�^Yv�c���ޏ,:�ǮS݁��V��7�V��������   `�3p X�.i4��*}�(b9u  ��T�!{��*#1zV��k�C���ع{_�Tw`��d������w|5u   �r� ��u�������צn  ֮��]�|p�q�1��c�����c��Tw`�)eY�n4~�kj��n   X�� ֠ˮj�5ى���ʞ��  X�^��r�Ygf��;Xy��C��c����N�b��1<��Z��m�3�[    �w �5f�ιs&f�n�t�H�  �g<���s?���`���<;��8�LN�<u���g��8#���K���   `91p XC67Z��MeE��n  !���P��s*>�唘�	������Na�� }}a�����=;���   `�0p X�X=�/�61]~k�  ��W�<2P�J�;X=ڝP��p�ܽ/�,,�"u���JY�q���[��S� ���f    IDAT   ,�  ��E���6����3S�   <�׽�<�3�j�V�x�h����}�X�ESw`.��������d��-    )� �b�w����d�͝^I�  �X��̬���Rw�������}E{�C���1u�����CՁ��}�Q�q�   �T� V�K�/\<1[�8/b%u  ��	巿�2������	ž�c��}yga!8�Xv��lnӺҖ��}+u   @
�  ��{�˧������ͩ[   �GV
�o��T������#�:�?�/oON�<u�O*��ކ���[vܚ�   `�� �"��c�v�f��n  8?�s��'�����`m�����[�����Lw`��J��n�������o'   `�0p X%.��u�x+~���6�n  8Q/8+�������m�͐�{޹g_��y��{ Bah��n�y�m�3�[    ���; �*�uW����v7�n  x"6���缾잆e��	ž�c��}yga!85Hn��׆�y�o��K�   ��� V���ߞ�ʶ�E��n  x�J�����h��5�G�!>t vt_ޞ�y�`m�V���u��=����   `1yQ  ��}dGs��d���:  `�;��塍�3�,ݻ~�����Lw �r)랶��n����O�   �X�  V�K��z�X�g�«R�   �*/}A����j�;�����������Cw �,qݺ싷7��N�   �� V�+n����//,�g�n  8�������.���Ќ�=��{��N����X{F�����W_��uR�    �J�  +��Oο|�H�s�NX��  �T�TB��WF�g׬ �N(�}���u_��t݁�5\�׻���>��   �T�  `������ǎ�]y�S�   ,����246*�;�D�y����ܓ���P��֎Z-;����ݗ�?u   ��`� �\�hn��>\�PJ�  ��^�R�9�(���+�:�߿�h��ECw`I�U�溑��on�q�   ��e� ���qG�����OL�ߚ�  `)�����//������{���L�S� �_V�����m77j7�n   8�  �Tco\�H����R�   ,�z-�~�-�=�fuȲ��;�.Z�&��;���R)��~kcy��F#�W$   �� �eh���s�&�?l���-   K�W~�2<X��p����;�)Z���^�`u*��_m�w[c�L�   �e� ��\֘{ۑپOu�q0u  @
�����ӟZ����29z?�'o?|0vS� ��@-���n�^ߗ�   �D� ,#�l}db2��(b%u  @*�~zV}�K��;`����Z-M��]�����N�   p�� ����h,�Bt�  �i�CY��<�����T������X�R�Y�.�yG��S�    �) ���X:��?31ޚ�  `����TFj�������;�XJ�,߰>�r�յ[S�    �4�  	m�zhp�:������R�   ,'oxUy�)��j�H��XY��F��zg��-    ���  �Fcn�C����lfOO�  ��<��Y�ϼ�\O�)��a�H��#/�}��fy�   �Gc� ��eW��o�?j���S�   ,G�ǲ��XN�ˁ�;p�e߯V��{[c�L�   ��� `�]v���M�>��C  �ǐ�Bx�[ʣ���sl�݁S�^������é[    ~R)u  �Zr�΅���|��  ���"����K��������W��y}y�􍡒�Xٚ��ss�?���R�    �$'�  ,���i���D�,���  `%x�sK�=�TK�����������T�S� +W__�_7ֽ�����N�   ��; ���Ȏ����y!D�_   ��I�e��_SJ��Y���������ٹX��V�r)�n\_�����R�    X ,�;�}�p�sS��M�[   V�r9d�~{e$�<ˆ�&���;��a�n���;p�J�,߰>�r�յ[S�    k��  �d��C�3}#_��/�,u  �J��7��֏e���R�E����?�'ow:!��V��T�c���?��vI�   `�2p XW�4��c����\�xz�  ����/.��zfVK�+M����wݗw���81�F�_yi�_=7�S�    k��; �)vō�<���	R�   �tO}r���W�Sw�J�j���{��}�N,R� +��`��ڿ�onkl�I�   �-�  ��Ǯm���D鳝^J�  �T�C���VFb�<N��|ȿww�z�@���k����o��x8u   �v�R  ��^�>��x��v  �S��qf�N��`(��g˃oyceh��Y%u�2,����ϗ���{f_��   X;�x p
l����ȱpa�B  �S�U/+ןuf֟�V�#���;���t�S� �_�/��\xsc�/R�    ���; �I�|u{Ǒ���k+  �E��3��_VH��M����ñ���f+�K	��*������e�4���   X݌�  N�EW�>9>�M�  ���ү�SI��U^�x�������v�b�`�*��޺u��[wԿ��   X�� ��F#��t[�75����  `-xǛ�#�ZVJ��Y��;��[�=;�y��c(��|�X~�m���S�    ���  '�;bߑ^����   K��D�n�ծ�J�xqy�-o�=鴬��X��"��'��?{w�&�Ux��{##2"��w���J[I���.�d6��v��{��=v����-Ƣ#���0�jl==��=m76[c�LӶ��AІ�c�ReefU���q�c�CI��������R�9�w�Wn����-   ��d�; ��p�M&�k>0=���  �������{Vl�����hZx�Kݹ�i�܁�o���_������   XY� ��w��������\89w  �j�vM(_uee(w�6)���3��ȗ�͹fJ�{�޳n8}bS��_��D/�    �; �Q��ߜ�v�@�ósiG�  ��(!��++�վP�n�ը��/=�����Nǜ;��m�����Hl�n   �?�  ?�on�2֊�o6Ӧ�-   �ٕ��6Ǿ����̅�#�i>�tZ�����������뮭3�[   ��ͦ ��;�_r�?d�   �C���V��z(/>�������kC���S3��#��{��i}�   `y�� �x�ms?v�p|o��[   aӆP����`���b鉧��Ïv���C���zzv�pzݝ77���   ,O6� |7���ԡ���n�  �w��n�-�Bܹ#V�����c-z���q������xs��-   ��� �\���t�p�v�[��  ��t;!�N���w�TBq�e��W�C�6�J� ��f�8:>|���9�[   ��ǀ; ����m�׏��[���a,  @:4ڹ��o�p,���%畍z��{��Za��T�?�鎹�s�    ˋw ��ߍ�̿m�H��]��   z��X׀;���Bܹ#V_�b��ݱݲ���������;���n   ��3  B��������gsw   ���UB��k*���6,33��G;s��K^N�U�,����[�{���n   z�  ��62�����{x����-   �W��Z;����;0��bgnv6ts� y�"t6�Kw�����n   z�  �������L��L/��  ��[;\����J������jY	ql"�S�],��f���kn����;ȝ   ��"w  @��`*7}�����xY�   ��C�v���+���.�_sU9�c��T`5�T��r��͛r�    �ˀ; ���}w�����?9</��  ��w�P0��X������W\X4�U�j�R���ŵ׍�ݒ�   �M.�U��S��O����tؗ�  �f����\��� ^��[b�k���9��EO�`UI�n?\���ߚ�   �=��U�=K��=����t8?w   /��x2�+@Y����X��������,����������:���-   @o��  ��/�;�gG����g�n  ��;��X��%e#w�xb�O����4�!���Ά���ｽ���   @o�� X�n�����h��  V������ ,��B�u\��������/w�t�������o��    z�w `E{�;Ӛ�r�M���s�   �x&�R�9��;���_�%�/��h4<˂�bl"��׿m���   @~.��Ƒ���͏Nυݹ[   X|c�wX��n�}���2��Բ=тUa�H�*C�   ��@ `E�qdb�t���3s��-   �&�����U!�=-�_uE9�q},s� �����U׾m�wsw    ���  ���͇g+�m��[   8v6����//�rw K#Ɛ��Tj}��Ns�R����޻����FFb7w   ��lp V����yb���  V��#���r��"�wk���2�kg�����ɩ��s��&_o   �Uƀ; �b��Lo}j��gs͸=w   �^�0v8�sw K����.��+���kŰ�MN�n�BӐ;   �2.� ���;�N��n6��-   ,��N+��<������^H�o�ҝ��c���8v���[��>2�]  �U�w `�����I�����   �ϡq�a5���x�Ye�e����^�RMN���f?42���[   �c�E ����;&O���k���[   Xz�㩓RH�;���l�}�yYeh��X��~��49]��lk����X��n   ���;  ��z�]S{������n   �W^Y\�&Trw �al"������T��n��`���������\�   �ذ� X����ҩ��  B�vr7 �cúXyՕ�ОS˚m��LOǳf�>d�;   �\6� ����>�kv��ps>m��  @~�o�}��_�� z����~���#��Ê3<��W��##���   X\�V  �ʵw̝0s$n  �=7��1����=����+ms�ir*�}v~�Cwߝ�r�    ��U �l��ι�s�Ň�[�p;   ��5��T�����"Ľ���+.��2w�x�g��?����_����6   � ��ead$m�:>�l�M�[   �=��S;w��֭	�W_Y<�̲�0
+��tط�����$Ͼ  `�p� z�M#S���m�i���n  �7��u;���c����_qy9�v�m�RLNƋF���7�   +�> ��F�J�U?:�L�s�   лF�lp����X�����S�Z��V������f/w   �⹲ z֍#k�m~dv.���  @o��	ݹf��� ��C�{Z����rphИ;�G�ʫ�}�����    ^�u @Oz�;Ӛ�f�O���	�[   X�[܁�m��XyՕ���]���x�&��+����۹;   �΀; �s��h~tv6���  ��cl;�e��U6^vq9P�����������|w�   ��qA ��_~w��7���'�n  `y98���n ��-�b߫_Z<~{����8���~�ۚ���   x�� =�ߝ곣͏N���r�   ���
�v;tsw �[��K�/.�W6��s� /�����ni�3w   ��p z�{>�j3�?25O��  ��!�H���b��X}Օ�ЖM���x��'�v���-�;   ��g� ���S���;���ٰ'w   ���xh�n V�F=W]R������e��n7�.ᆑ��s�    Gǀ; ���w��������tyv���#!�vr����r�  �-��;6��*�w�k���Z�6��{��/u�qt��7׏̾!w   𣹄 �y�S9���?�����nx>֯��VN<����R��?�m7�C�� @���=cwQ�1X�,�Z5'�,�E��xj;²��«_{s����?w   ��p �IEw�'�ⅹ[ �V��9{�����z�穢q����Գ��n�.  ��m�}�z�S`������}KQ98�m�Z��a��͹x�U?������·s�    ߟ~  ��v��''�E�; �F,Bص3V_{Ueh����wnm�cq��@�b ��0:�zS�ք�+//�N8.��n��nJ��X���o����-   ��g� Xr�����#�չ; �ƚ�X\z~�qꮢ�,�s���5�����ia)�  �^�2��;�j�`e+���VT�cq`4����E��J)����W��-O~����w�{   ����3  ���o�������; ~��qϩE팓�Z�Gv�£i�+�贎e  ?\_%ğ��2܁Kdf&t>�p{v�p��n�^���k�/�������   ��"w  �z�8Ҽ�����; ~��Ǿ�^]��]�?���B8{O�o�+Ǫ �m�ґ�d�2�dB���+����,�N�:R����1{a�   �[\� K����~��D�>�d{г����|_ٸ��r����Fb���Р� ������c�g�Q�_zQ9P���`�h�S}t��?�r�Ԟ�-   �7�\ ���>�3�cŻR7��[ ��X�p�	�z�e�,�43:yo{��
i1�<  ����}�[�� V��V�>�����%/��2Q����5�����c�[   `��Q 8��8�|��X���@�Z�&����2x�Yec���C����/=�l�� ���C6��Ԫ���r���e�p+�B���N�?I�s�   �jg� 8f�����;~��M��- ߭,C�{F���+*��քʱ�ol����S��? �n���\3trw �WJ!�>1�^qyeph��ϰ4�q��s���L�   -�vB �o�+�<}l����B���ݶl��}{�����|]�s�tf��xj-� �o����q�k �N'��}�3�ؓΆ�6���~rd$�;   � ,��9�s|��~��@���B��ܲ~�%��R���yg���룏� ,�C��v������.��W6*���Mφ3�����uL�s    � ���idj�ԡ���VX����������2��XKii�	b�ʁF� `)���@Oٹ#V_����5K��5��LM��7=����   ��  ͛ޙ�L��>�lŭ�[ �A�?W^T\xv٨��;��Bqžr�,m� X*�3��j�n��o7P�+���>1Vs� ?��#饯���[�;   `�1� ,��|,�Ə�hz�{B��B�E�w��k��m��r�����X^r^Y�Nb  K"uC84�:�; �[�!���l\r^��"4����᧮�u���   ����! ��y`���3���- !�04��/(v�PԊ���cR�R;w �jШ�b릢'^x�nk�c�s[���x�3?R����o�{�z�[j��s�s�   �j`� xQFFR�}v�&���- �a���z����`#��yg˦XNͤ����� ���p�΢����VCq��Euf�9zVJq�/�ꚛ������  ����  ,o�:�39U\��`h0?vi9x�Ye�챭��-���]6֭��1 ��6v8u:][���V�!^|n9p�e�pR���R�c��o�e���n  ��΀; ��]ws��#�U�;��-!�9��]�rhúX��s��"����������  �]�0>ڹ; �Ʈ�b��W�=Ã^�����*~���|y�   X�\� /�#s�:>]�Td�~m,_uE9���X�����?�z,.���� ��z�`��-���v8T^~yep����7�&�N��M�����f��n  ��j��  �]���4>^��M��r@���e�Sc�rl�nO<�Z�=ܙ�� ��5�8�欄�:P^1z^�!}������v溝�5�w�V�������_���)�J    IDAT   V�e? ,�7�4_��H���N����N�á���J}�pXQ��𷝹�|=���  X6����՝�c_��K�@o�H�O?ԙ�k�n��;�������k�:��   V� �Q�qd������������>�ᴓb�%��+bk����}�3�́�� �Z�e�6���+��o�}+�w&��Z�{�:���sf�^Ө�ǆ����7��r�   �J� 8*׍�7=]���VZ��X}�Cq�9ecú�����v;t�����ɩd+ ���B<aG��:����e���#=�����W;�N��[���[�՟��v  �"pI �HozgZ39����|ؒ�X]b��c��}�����2*��o**�?�]�tr�  �.�Nc���'R�݅n7���X��E1@ψ�7ľ�kc�4���w̷¶P���'��X�   X	\� ?��w���=6�gӳaO�`uŅgW�6���-K��XZ��}��  �*����N�YV7o��ܩ�af&t�y�=;9��Cټ6��o�^�-w   ,w.���n���#���;����b�{�z���-�|�����_����  ���P�x\�w��Pk����
�N'���Й}�ٴ����Cڸ1���V���-   ��p ~�ko�}����'rw �G�?��)[7�U����y苝ٯ?�Z�;  ��X��}K��}BQݶ9��dcH_�Jw�ѯv����(b{�t�]�����-   �\�x ��n�����K�;��c��X�wv�语ޭ��-��>yg����� ��j4Bq�	Eu�΢Z���s`4-|���l�R� ��J�۶�������s�   �rd� �7����C��nJ��\Y�xΞ���]�j���j-����mOOM��  zTQ�p���w�β�yc���bf.t�y�=;9:�[�j�xx`M����m��r�   �r� ����������tS_�`�۸>��W6����ˎL���?ݙn�m� �uk�b�kgQ=yg�V*��K��	��/tf�z6-�nB�����o����x�   XN� ��;�_rp,�I��[��-!�����uj�ѹ�h<�\Z����L�� `Y諄�kg��zbY�B'�tb�ѯv���n������Q������   ˅Ku  ��u#���,>���s� +��`(���8�X3�~�c�J��-  �h�nc���'��C��_�qh0���؋�����u�|�`jw:�s`u[h�������ù[   `�p� ��FƆgg�k��r� +ۮ��z�޲^�"/D�!}����O��< �r4<�SN,j�vƪ���R���O=؞=|$s��֯����o��   ˁt X��;�=�x�O�f♹[����㾳�ƶͱ/w�r���W��L�N�  ��j5ēv�ꩻ�Z�?�{�����/tf�|��ҐS,��a��;�y{��s�   @�3� �������������ʵuS�\tn���;��9�yO{z���[  x�2��ž�O.kk�C%w�r�җ�ҝ���fr��lbi��t�{n��A�   �e�`��m��=q��������:��߳��g�E7~8���3��N'�N `l�*g�.k�6�JJ~?��3R�w�:��0	��Eloߔ�{�[��[�   �U.�`�����M��ŵ���{ Xt���伲�~m���z����Ý��  ,��X�rbQ;��X��>���L��=vffg}r��3[7-��w�y��-   Ћ\��*t���O:\���Me�`�ٹ#��{IY�TB��e5��/w���ki>w  �����]�v�	�V���E՜�{�̌M�N�X��kql�@����x0w   ��� �ʼ��{���`���[���,C<gOٿ��X�ݲ��ҧ��>�?-�n `��UB<��X=��_�)�xR
避I��?�q��L���k��׌��V�   �%���*2rW�x�P�p���nV��byե����b_�U(��R�={��n·�; ����ph<t��x�o�bwx(�}6�� ����B
qt"��(a��a}�l_�Ч��H�   �%.�`�x��R��O�lj.���X9b�i'��KN/�ct��i�:qO{zސ; ��V�!��#V��]�,����S��w�:gJ�a����u{��   �+� �*�u��&���;���V�s��[�{��XX����3��� �c-!����<��_;�/�đ������f2�K,Ɛ�lH�������   ���; ���2�����_�� V���cy�y�@���-|��=��?�Hg.w  K�[��em�p������|���`gfl"ur��jS)bk���~���{s�   @n�`�����������}�ŋE��k/9����Wz�翔f���N+w  K'!l���2��H�nH��3�Գi!w�6�jqdpM�����c�[    ') �����K����	��-��W��xɹec˦ؗ��.��3s`4�s�  ���n����(��/T�!=����#_�6s��jS��n\_��]o�Gr�   @.�`�����Iͩ�g�a(w��m\�K�+�X�n��B���v���S7w  y|sн���e�`yzzj����\�R�XM�_�^����Ht�  ���R V��FƆ��ji·��[��-!�~r�]|n٨�n_N�2�m����Ow�� �J�3����R��d��e�oz�����M���`Xh�F,�V+nI��	|�?��   9p�fd$�����xJ�`y��B���r���Z����U��X�&�O�Ov� �R)������S�55�:��e�/t�Z�?�o/����|���J�U�v�5o	����s�   �Rs� +�X���tyv�`yۼ1T^���ЖM�/w/ζͱ�%����;  �+uCx���_��=��;�s��;?�Qk�Cy��������,X"�ۍc��7�6���-   ��la���7�p�P�>w������Y�mm_9b�ϧ�ǟ�,�n �7e'�ս���ժe8���tC���������%,��J�۴!����Z�b�   X*V `��ad�'��f�&[�����E��[c5w�/����3��C㩓� ��Q��x�Ieu���_�� G%}��N�￑�s��jQ������52t0w   ,�� ����{�?W�@��[��i�P,.��^�Y������mO�Άn�  zK�?�=���O����p��x����\r%1�H_����ڑ����   ǚ� X�F�J�
j-���[�����˾+.,�k���±U���ecQ>�tw!��5  ��v;��S���i��㚡X����~m����3ϥ�3&{����]i��Ч��g�[   �Xs9 ���H�>;7��鹰;w���"���(�O;)��nai=�lj}�s���  ����cyΞ��a]��nz��Dj��`g�5���ذ>��{G���   �cɆF X���`�x!�P���r�p��t��X�sjY�� @�:4�:��3��:3�s����]��ʫ�����161Q��u�L���   p,�� ��u#s������X~�l��K�+��^W�C��������B�  z[Q�p��X�{Z�_�s� ���B�~�����C���V�JZ[7t�կ�ܸ/w   �`���kL��t����,���S�ڙ����,@��	��nO>b#'  ?Z���e��]��3�ݐ>����a)Ԫal���5w���   ��4 ,3o��y��\�hk!�n��J%ċ�-�;��j�z��\�~����\3��-  ,�C�x��E�����?�i��7�|�X��o'Ϋ���hy   +��� ����LO�����Vڐ�X>�cq�%�����/w���/ƍ�c��gRˈ;  Gc�ғϦ��é�nM,�k������ms����sc��5�i-�M�&;'<��;�<w   ,&� ���|��hf&���X>vl���^T������@�z,�x��O� p��gB��O���\�n�P�e髱��l\+C�x湴`���f�8�W�u��O��P�   X,.�`���ֹ;'&����Xb����KN��)�����£i�+��rw  ��Tk!�=���}b���o��`Z��C��Nǘ;+�"�6n����on|&w   ,�� �\?2����;�)��7�#U*!^|nY߱5Vs���O�י90�ڹC  X�֯���{��������c�}���Vː;+�j?a��ꑑx0w   �X��ǽ宩=�<[�H���[��7<��/(�c�����ݿ�Tgzj:us�  �<�"���c��g�z��>Baj:u>qgfv68o�12�H_�`W�k~��B�   x1� @�ndlxb����BZ���};���K/,�u$�pE���E��g��N�  ��������b��2Fw`��Uc�s{Q�?���6��1��7L/tNz��w|,w   ���G���b�U|`f.�����X�p֩E����zQDC#�h�j(֭��Ϧ#  �P�n��S���ڡ�hx&�]_%;�}�R{���	�B�U�r�5om���;��   /�͎ У���>9��������s�ƙ��)و��ٺ)��}Fٟ� ��or*u�����әm�B7w�W���/+�m���-��n7NL��x��e�[   ��2  =�������xz�aU��i4BqžJc�p�@�c�/vf��Dj��  `e��B�{j�ʮXu��[J!�����Ϥ��-�U�ő���k�;�x:w   <_.���\�k3�O����I��-@�ڸ>���+jU_e��J)���Lg��x��n `�ؼ1T.�[ևc���*}�K���=��j8��k�T��1z�  �e��1 ����cr���}h-���-@�:���������v��Cܱ��{rwaa!��=  �3����'S��Iiӆ�RDy`��;��X�x�Pj玁����Z�����O�   x>�@�I��l���\ؕ��M�a��E��{�F4����!n�+�?��w  K
��x�<�lwax0����*7���Z5��R۫հ�����~�[;��r�   �Ѳ� z�hwf���@o꫄xžr`��?w����X^r^Y�N�  ,�����}�����fZ�����qʮ�v�9e��,���Ʊ���7�6�c�[   �h�� =�������Xqsɿ���������A���ѯt�_��n3w  +S��9{��]��Z� ��i���3��U��0�fs���~s���-   ���������a�����[7��e��J�ח�1���:�O=�r�  �rm�+��-��U��xj���L�L��"��o���zd$�r�   �c$ dt��������i0w�{N>!V/9�l���vzJܾ�����n�4  �ؘ�	ݯ?�Ze��u����Ҩ�b��Xy�ٴ��殁�c��u*�=~�����   ~� ���H*���΅r� �%!�=��?����!zOCܶ9�=�lh�۹k  X�R
��hj�v6�+�j�˿��4�ض��<}����䮁��ي']��_M����s�   ��2 2�οcr*�����������ƞ�E��a�X\��(K�`  pl������ә��o�f�"����P���r��>aML����w�^��   ~�A ����l^��h|_��|M�G��P\yQ��v8Tr���z�Ժ���l�  V��kCy��ec�pt����L���}������+Eݴ���w�9��   ��0 ,�k�;ab���N���G�ք�e���C��4X^�ǲ�Iil"�`<  ��\3�Ǟ���a�X�|`U�VCq��ط�`Zh�|�C�B�^�Ч��@�   �n�g `	��>���\+l����[b��}�`���-�Bl�TTO��ԴMz  {)�p`4��;��[6�j58K�*���q�b��Ѱ0o��|+l����6��ĝ���   �Υ/ ,�-�̽gz.����ݻb��ˁJ_�u��,^|n��  K��x���Ov������+���X\}i9�n�%^�X����M�X�   �v�h `��xG��L������X�pޙe}�������L����i�� `�m�*�[����j�n��'���O��-�T+ar���5w��x&w   �`� ��Ϳ9�SO����N��-@~�J��]P6�n�}�[`�K���3���K  Xm�2�s�����Ք<�������=vfF�B;w���v��_32��   ��M& p���c���/-|x�6�n��B|�������Y�������`2`  ��J)��S{�p�l�XT*Ce�;w}�GRgz&ȅia!nL������[   ��  +ݗ?3�{s�x\� ���X�����������Sv�ݻb5w  �ӳϥ�_�ә:0�r� �VY�xžr`�w-�O�����g~*w   �^ ��#�׏���rw �m\�+��ժ�LYR
��wf��� �|v��������<V��B���:�O��b�X�J���?�w�5w   ��] 8F��k3��}����d�-�r�o�}�[6
�2����O��gg}* �|�Cq�e�״`e3������_{��Hl�n  `u*s �Jt���ڱ#�-��P� ��w�څg�����T��n��ǟI]#�  d�j���ө�6��e��V�C<~[�wd*u'��h/��BX��k���=w���-   �NE�  X��[�ߛo��;�|b��3����(�)�`�Z3�K�+�� ��R7�G��m��g�3s�d�V�C�����c�/6��ux���Ʒ��Ϲ;   X�� �"���[N���ȧ,c��ܢqܶX����o��m>��n3w  T�!�{IYwf��+��>������B�X��2�o����w�y��-   �.�`�q���g��I�T�n��B|�����6������O>c�  �ްkg�^����g%�r���ߟ�h̾�#&s�   �z�H< ,���魣S�7���U��������{��E甍�' �	�=�Z��������,�C����qܶؗ���f3ni���>w   ��� X��`*�Ni6Î�-@k�bq�e�����]�Abq�����g��vH�{  `~>�ǞJվ��+O�!���;2���ӡ������x�+^{s�ٿ�㳹[   Xlp�E��K�	��� �ظ>�W_Z������#��Bq���Q�1w
  �B�tB��#���>ܙi���J���w��/��x���n��$w   ��� x�����W>=��?�^�Ui��X���r�,������gR�wfsw  ���ť�k�}�V��B����̳ϥv�X����P�1s�{G6L�n  `esA /��H���T�۝T��,�];c����FQn��k�p,;ݔ��N�  ��VH�?Zվׯ���=��1ĝۋ��S�;5�k�B�ۡQ���=w~4w   +�M� �"h��n��]��Xz���)�1n��=e�O� �k:�>�Hg��v�!��O�!^v~�p���dq�u#����  ��f� ^�F�n��.���,�X�pΙe��g����Ë�R���[6֮�u1  z�cO����mOOO���$�0�m��4�u�Hy�[�ړ�  ��ˀ; � 7�>{�����sw K+!\tvY?�؟�V����+�Z�#  ���GB�/>՞~�����,�C���r`�&C��Bt:�66Z����N��   �1aK <O�����O�?n-���-��)����8n[��n������kc��3i!��5  ���ڟf���msQ��˙�����Eߡ�ngf6ts��r�j�����	~�?��  ��c�; <O_�J��fwK����    IDAT`�T*!���Jc�h##�7ľ��,�;  �y������t�g�AXX!�"�+.(֯�^������m�u�;   Xy���p�����ɩty�`�Tk!^}ie`ӆ`����'�ک�J_I  �g�M��_~�3up,-�nG�/Ɨ^\6��_��G�[�z���%   �,��(��ߥS'���� �N�?W_R�[*�[`�8��X߲)�; @���ػ�0��¾��{έ�V���[��ZB-�]�Z�Rk��x��!c3��8����lbp��16q����d&�<��䟙	�m�1�M,a!H�Q���ֽU�ު{�;(���VW��n}>����|���{������!}���Ï�^�!��^��P��`cz˦��)��A�9܉�zv6��  �	�$ 8
�~_*�Gz�����nN�M3�x����M��of8�bq�E�Ciue�X �!�B8t8S}��XQ��;	xie�g�cO|'�����c��OS�M���?��  �h�5 �_X����x^���ؼ9����1Ӝ�B(�0>�����c#!  ����N�򑪽���-�K75�:ؘ������B�s�Ͷ_��  ���� ��_�{�ϵ˟��������1=9�2�43ʃ�ʦ�� 0�Z�T�ч�o?�Vs� /]s*��\WNOLx��E�S�ꌽ��w�-�[   X��H	 /`v���ۋc����d�`흱-6n���k��0�4˲��;�� w  �����N�u�iǶ��0ֳɉX��-�}�PZ�|��ZU�f�=���=�%w   뛁; <���T<�K���g�n�ޮ�q����tQ!�0�vZ,�K�n-�:w  ����#�j�S�sG1VDח��MN���b�O���)�^?�z叾�����d�   �/'S��8����.����sώc�.��� �NJ!^��l�~j�6  �·�L��o�Y�&�XX�N�7h4��-#8s���|g��   �_� ��t����ksw k�e�ʱ�2n�ac�7\SN7��a X�[���T��� w��l;-��t��.�vG�����s�{��i"w   �[1 �n��ߺЙ��Wi&w��.8/��S4C0n�a�h�x��E����Քr�  ����{2��L�b�f_$��l�˭�b�Ci5�&��2�MˇWw���{ߟ�  ����w �z��������ںhw9~��TJ��^l���-�rw  �Ѫ�>�@���/W��ba=;kG�vO9=]��6�*��7�.�&w   �[0 �=n������xm�`m]za9����4n��g��8~酥�[ ��|����������`];��8��r2w�).�˷�~v���%   �/� �����/�k���� �֥�W\� �ؕ�ɳόc�;  �X<��4���U��n�r� ���q�����(����~����   �/� Bx��R�����JL���bҸֿ�B��uK(s�  ��X\�}d�yz.r� �o���������^t��%���g�   �w !l�Rﮥnܝ�X���ˋ�K.(|BFDY�x��rzj2��-  p,V�!}�u�[O���-��I)�}W�Sg툍�-�^i�x�����   �� lx�r��u�V�wrw k#!\se9���
_h�Ӝ�������9�  �3U�����z���R����������#w8
u����տx�{�X�   ��  ��l?�I�au5m���x��+ʩ��D�vQͩX�L���Ci5w  ��SO��r/��ۋF��׉`��1�];��w�N�n��*�b����Z�������-   7'��������;�ϸ6�s�.�/�]���  ����ci�C�,���:wp�c1�t�1=3�+�����n�m�"w   �͍ 6�;޶�����;�ϸ6���ũۢ�� �.=�t|ྪ��U���MN��6��&�/1����T�:c�~׿Mӹ[   ^� lH���o}�]ޓ�O?è1n�+�pM��4]� �.�;���}Uga1r� Ǯ9ʛ�-������W�i�}����;   ^��!�V'~e%���8���ack4Bqˁrz|ܘ  ����K���N��[�c�ush�rm9]�.K���-�����+w   �����wu���8��8��ہB�����ʦs� X��*��_-}�������O���*\�J���x��o��s�   0|�� p2�~v������4��8q�ہ�5ӌe�á�i��  �K
�Ci�BLg��r� �f�XNM���w\����4Y���O}�����  ����  6��J����4��8qb�5W����q��s��  X��j�����B�����ĉ�/,&sw��[X�׾��/��   `���a�av��N��2wp��"�k��ݻ�ہg�wE9u��ї�  X׾�XZ��g��6r��沋��^��kx1��x�/��v��   `x��!�ڻӅ���� N�X�p��Թg�)�o�_N7��} X߾�dZ���W���P�n��՗�S;ψ��0�Vi����  ���!? #���K��zﭪ��g!{/)�v���v��M�����tY���  ^���R������d��H�!^���>uk��1x��pɭo�ߙ�  ��`����������x^����{Y9y��¸8*[7�����Tt �:���|��,-�*wp��2ě4|a^đv���ͮ���  @~n� 0��k���bxu����si9y��8��X_���/���w  ���r�?��������a���+�-���}a�O]���r�/���4��  ���Y���41߉��j�~�Qq�%�������򋋉sώ� ��u{)}�U�𑰚�8z�fby��r�p��W�w=�x���   �e�����Ǘ�ۋg�� N��/��:}x	R
q���y�/� ��!��'��'����a9��ظnoٌ����oǿ}�l��;   �ǭ F��������Gsw '��ĉ=��S�;���,B�q9=5} �u��R�����cO���-��۵3�_�r9��Iu*��u���s�   ���; #�;M�:q6�`�#����񽗖�'Ls*7�/���O  ֿT����Uˏ|���n����ύ�;`X��q{wr˻rw   ���; #�;��=�~:-w��]�8~͕�V��ԭ����!  	��3�ݯ|-�r� G'�����ڱ=6r���j���ݽ��  ��g��Hy�l��:��N���]a����Ύ�'rw  ������ރ�n�����הӧl	e�FuJEk1�����R   ���02�����r�cXX��<#6���l���3���^ZN���iy  ����Z�?���cH�[�W�!�|mc�����K����wߙ�  ��ˍ FFf뻺�pz��ٱ-6n�_N�h������M��1  #��G��O?Xu��a}�������q��๴˟����+sw   p�x��H����+���� ^��O�����I�h�����  ��G��V>�����;�[6���}e����luJ�b���{���  ��Q� ��jv6�j��j7�n��)[B�CӍ��0��o|<���ǞH��?  ���V����>{G��0�f�������Ci����`g�W;���=��  ��g<��w8���[�;rw �o�L,n�ָ�k�iql�%�T�  8���j�����S�*'��wŉ�ΏN���0ߎ��{����  ��3 `]��{�7�Z��� �_��W\W�LN�m
�w��b���x�  8��vZ��g��a��{i9������&թ\l��z�{�X�   �V�;  ���l�3����as���LM����3����R`h���h<=����P�n ���	�|+U��,�b1w����;��'����S�{������O�����  ���L ֭#u���^<3wp|��C���bff�K��p�1ăW��f�53  �����}�����ï,C��@�91��A�����6��7w   k��z ֥_�g���b��;��S�!�rm9�u��ہ�41����Ӎ�!  ���֏��P޴��.�A��Sթ���M�   #� �Ϋߗ�#��ݩv�3�GE�M���[c#w�ٺ9��.�ѕ3  #��֏�N��W��0l���ˎ�ޯ��   `mxL������{���+wp�b+����X�����8v�E�d�  8ў�N|��F��{v1~��q"w��V�w�ۿ2w   '��; ��ޱ����v���콤�:��b<w������Ĺg{1 ����!#wX/�^ZN�u�kS�^u��Z��{fg��  ��q���������0�;u��[�cw��ą�'M�NJ!�S6O;%��[  �D3r�u#��ln�\���X�����ʛrw   pb��n����ot����;�cw�9q�ʋ�d���U!޸����t ��y�P|���rF�0��2ě�7�!�n�a2ߎ���ޝ.��  ����< ��տ��~:wp��>3��SN�����MN����e�,�u ���֓i���_s*�7�/����0��#�{�"w   '��; Cov6O?��S�i,wpl���.�!���ԭ�q`O���  k�O��O}���h���Sb����M�{u��E���n��  ��a��Л�7w�����9eK(o>�h�q;0Z�9+�_|A���  k�����_�z�;�v�مkS�s������y�;   x��j���w�|�������4���mL7~o�i�%���3b#w  ������_�j��� ^�kS�~�*L��=�;   x�� j���wU�XG&&B��@czr�oM`������[��2w  ��/>\���hr�;�x�겹i&���b'�������  �K�f C�{���,{rw G�,C��@9==m�	��g��k4'&B��  k��_�z�u#wf�F(n�_N�5\��_�[���6;�5w   �����t�;Ӗ�BxS����"��W�S�n�Yd`㘚��Mg� 0�x��}�����<���P^{U9����2����;sw   p��� `(--��������՗Sg��; N�m����/+�rw  �ZHu��|�}��i%w�����/������b�����fۯ��  ��1p`��yO�ƅVxU���]za9q��
Ѐ낗ŉ�+�� �HJu�Z���i5w����8N����!�ꔊNw��W�/��[   8v� �W�/�O��;j�F��q��q�ʋ�d����^���fH  �h��>r�<���[��R��]U67�D��!���Mg�|�wg�   ��� ������n7�����Ƶ{�fJ!�n�-���gH  �說�>|���*w���P�pM1�h�_!�0�*�M��{y�   ���� �_���>�N�K���l�ʛ�7�1zX���Bq��rz̐  ����g�,-wS��xn[6����r*w�AUO�����;   86� ��~���D���MM���t���$���	��}e�9�  ����P�u����aH���/� ��!��N���{V~6w   G��v ������b'������F��\[N7�L7�ϙ��ؕ���;  `��;���'K�Քr� �m�%���3b#w�����_?{ds�   ��Q ٽ~�����Wrw /.!�W6�l�e��aw�q�e�ʱ�  �V�B����K)#wN�ڽe���LVV��PO�=w   G�� �K���+ik�����:s{4�8
)�x`Ol�~���  ]���'?W-�h��h|<7�/��2��-���b��;�Z>��  �g�@Vo�k���V��������8q�9q"w�zc�7\SN;- �Q���i�_I���s۲9���-�rw@nu��ť�;gg��4   C΅ ټ�}����w��=��w֙ql�%�d���hr"7�o4�� �({�U��o����s۵3�_t��+�ӭϝ�Wޔ�  �fP@6;\��n/�����S�����e3�L��ush8- �Q��/��'����s�sI9�������ͷ����{����   �����?��{�\'�l���MM���tY��T�v��K/,�� ��Ju�l�<���[�g�1���5�S�ѽ>6�A�&�����   <?w �t��TU0��!6��k���	�N�+/��g��rw  �Z������R����-��M����}�ttǏn�S\������   ๹u�I�ƻ�?��)��� �_,B8��ln���- �$����ln���
 ��ZY	���WK�~�s� �v���q�ˋ����b���w��4��  �g3p�z����ů�� ^ؾ+ʩ3�;a`-�e�7�/�} �Q����_-UuH�[�g���bb�����9���S����sw   �l� �T��z��Jښ�x~�'�?'N�� eͩX�pM1]8� �6�����Z
���MJ!��l6����-��_��w,���  ��s��������v��;��w�������N��N��}��S�;  `-=q(>�媗�x���P�xM���k6�T�rn�|G�   ���; '�r���T��aHm���.�!���`��}N��hw9��  ��WI�G����;�g;eKh�āll�n��ַu>w   �e��Iq���?�Y��� ���D�7][N7~�l{.�S;��F�  XK�~��:�Vsw �v��8�kg��9��[�|gڒ�  �g0����;i��o��<�X�p�Uesz� r�1��)��f�kt  FV�C�ا��V;U�[��R��,��f<;f�ZYM������   <�M
 ��`�w%���xn��(����&���P�r��1w  ���AH�}�Zꯄ:w��c1ް��.Kץl\��So~W���   ���~������rw ���s����ĉ� �0=����M� 0�:K�����R]����~[6��������K]�Ƒ���   ��Ǝ<�}WU''C��~zh컢����w�qz�s�1  ���|���|���;���ĉ��*��g�j/�+�xW�grw   lt� ���f���R�qe���6̈́�}�f�>90l.�'�?7���  �����i�ˏ�~��ٮ�267oe�ȥ�.~��ޟ|�   #w ���l_\*ޜ��x��X#ě�7����V��(�N?5  0Ҿ��ġ����~e���f��p6�^?���'{o��  ��5�&��[z��=w��b��ה͙'0�C�q9�l�n `t�:�O>Pu۝T�n��n��ґ�4x�u�S_��?�@�\��rwA.�V�����;?w  �F�{ N�_��{��⏫��a�카����8���������Wu�ʨ  ��53�W�ؘ�989�P/vR=���V]ͷR�j�*չ�`�l���_�|M�  ������u����������۵3��pM�L�o@���Ci壟��  e�O�W\ט��}8�z�P/,�j�����T�OU�\a�Q�E���V��7����n  �h�$��z�ݽ����!$���ٲ)����T�~��G_�j�~�᪟�  �҅���U��S�;`�J�N��Z��_����PͷR���"���P{����5���  ��4r 0:^��T.~�wW���o���6nX�.�(N��b���i5w  ���>��[6�b��8���YU��^
�b;��u5���#�qPU��p���i�·zw�ޞ�  `#1r���u����s��� �+!�r��>c[���KS�!}�Ag�� ��*�~��r�ԭ�!MB评za1U�Zh���B�:˩Nu�2�8e��:���{��D�  �����bv����ű?�O��{Y9y��8���c����W��G�]N    IDAT��X>  F��d�?zs�ir"�[�d����ϵR5���V;U�N0e�!�uK��߿{��rw   l� ��{K��\h�[rw ߵkg�ᚲ���| �dn!��cuǧ� e�N�:ؘ��}FR�tB=�JU���v]�K�~?�Ѓ!cH�NY�������-   ��� �d�߳|�S����NɉJ0$N����1S~���ǞH+��l���  �҅���U���ɺV�!�;�Zl�z~���Rud>TUe��Ms2}����+fg�/+   ��F�  ֿ�N�v�v!�t��4n]���[�z�k���  ��WM�S���g�[�hVSZ\
��B��Zu5�JU��d
#a�ϙo�_B���[   F�� /ɭw��p��p{��������X� �\��S���� w  �����Gn,g�nvhå���b��Z��_HU���v'��Èo�����y��8��  `��p��|g���]���-�3������b2w '�`�?���,�� �蚙ūnǰ�_�$��鄺�IU�����T��n/��a@�lN��W�L�.w  �(3p฽�7z�{d>����3�<#6n>PN�� 6���P��}���J0�  `d���\�k+����B=�J��b]�=3f�����]��9g���;���P�  �Q�s� �_��{n�H����3f�Cq�Ue3x���LO��k��>Q-9� �Qu�4���u���|��ce5���j-�j�����Z\J��*�Ť:�ss�=!����  `T@p\~������ă�;��2����ٺ�ˋ �W��|����  ���n���>��8������f�>�J�b;U�v�[�P��+Eڹ��'���-   ����cv�]�)�}�R��ẫʩsώ�; ��3Vˏ|#���  ��2>��TnjNE�&y.��	u���V'���:2�^J�À�35��՜�yv6z]  �s�' Ǭ��2n��p�9qܸ��t����bgP?�t�n �����㟭�^y}9���6��BZZ
�\+U�u5�̘���`���^<{~S��C��  `Ը��1���k�z*ݛ��ԭ���3E�7 ��_	�d�Y^N `d]za9q�Eq*w'�`5�ťP�-�j�UW��P�/���r���x\8-���ۿ�c)w  �(q�; G��Mc��Z�6�GA~�!޸��4n�M�������>Zu' 0���H�?mk��yF����za1U�v�Z�o=�Wx�!�_I[��l���[r�   ��( �ڭ��7���8wlt�����m����8�V>��j� �Q5>��Ҙ��e��K��B�j�z�����T��n/yQXW�2��9�~彿�|"w  ��p�; Ge�wҩ_����@����0n�Ŝ�#�_~QQ?�店�  ���JH�L����˙�4�R
ii)<3d_����T�-��W��QPUab���
!�|�  �Qa��Qyz�{��j1��6���e��� �����Xl����j�  XOϥ�sU��.+�r���� ����o�j~1U�T�ڡ�u)`�-.5^q�o-]��_��l�  �Q`������?,8L�������e3'�ptR
�����Y�:G�S��  ��WM��R���xw����nwB�j�z�U�V]��;_�-��S�[   F�q /����ϭN�&wld��ו��O��c����?<�t{�� ��4>��TnjN�"w˨��C�����V��Rud>���T������|v����  �������'�&��������.,&sw �~�-���~��T��	  �i���C���$����B=�J��b]�-�jn!T��O|�������䍳��!   /A#w  í�T�%��!��m�qم�D� ַS��Ɓ=E�㟭�s�  �Zx��0��#u��p��*�V��{�SW��T��/��n/�o�_B���[   �3�E �׭o����#�-�;`#����Go.7MN���������WI��  �b�+�3����z�P�;�j�S=ת��V�Z�P%g�P��E�+Ǯ�ߍK�[   �+7� xN��i��v�u�;`#�E�]]4��8��^ZN�����o���-  p��:��?P-��͍��{O����b��Z��_HՑ�0���c�N���z�c�k���-   ��xN������/.wldW^RL��6 k��B��G��V�r�  �Zص3�]����ݱ�R
ii)�s�T�/���b��Z�Z�cv��E\�|Z�c��-S_��  �9��g��Mۿ����d�c{l\��b¹Z ��������}h�Y�� ���֓i���{W���r�TUH�v�Z�P-��zn!UG�㠪��6�:��+�l�aR   ����g9\��]ĩ��QMM�x�Ue3%_�`�LO�r�9��ÏV+�[  `-|������Fcf&��[�U���b��ۡ�_���V�:˩N��/�����b���{����_o~,w  �zc�����+?T�҃�#!�[4'�C����w�9a��G��;  #��B�����X��8�	���^XL�\+U��:2��n/<k���R�T,-ŷ�~<w  �zc���i-��-�iݝh��ʉ��X� 6�-�by�)�<2���-  ��R��_��e�+S��V���ja1T�T��NU�x�o]�[������  ���i �|w�ӽ�[O�.�����Sb��7��b ���?���?Pusw  �Z�E�<XΜ~j<i?UUH�P-�S=�XWs�:2Ue���LM�'w5'o�����  p�����0�o5n�<��+��� �l���<z��F 0�R�������Ʀ�<��^�P/vR=���V]ͷR�j�*=k��'7�F��ŝsӽ�!���-   � !�n�]������������殝q<w �g���FZ��  ki��q|��e�����^XL�\+U��j�S��'���&'���5������*w  �z�w B!,���s7�F���8n�@N��)����� ����cie���8k�Q݇I�N��Z�juB�خ��si��;��c��mg=�}�=�[   �'�n�g�g�z��;wlD�7��Go.7���e ��M�CQ����� }!��-�M�������CjwB��N��b]�-���|��ʘ�g|�h��s�߽=vs�   ;'�lp�����B�'_Q�p��i�@++�~������~U��  �1��!}�s��mEc�UW�P��R���e ����zKZX�#���)  �aL������7n����ˋ���WL�� `cYY�Ï���_�V�H	   p򌍅��&���_���-   ��	� ��l���{�;`#:kGl\��Of� �$��3���|�Z�   N���0����g!�_��  0̊� �3z��_	��fj2��{�fJ���ګꐾ���?8h��o�   ��B;��7��ҙ�;   ���;�����[������=Esb��0 �\����_?8h�����b�   �[U��֑�-�;   ��a���G�oY�����\x^9~��8����v�pZ��U�����^�s�    �]���U�8�۝�  `X5r p��1���T+�����l��ŕ�ĩ� ����4�����SO�A�    �[]��b��B�{�[   ���6�~=��A&sw�FR�!\��l�e��[ =�v�>r����T�v   ����7�qo���   ��	� ̭��3(�h)w
l(W\TNn�� '��j���H����Ou�    �V]����Bxu�  �a�w�f�	w�4��6�m�����ǉ� �����GS�������G��   ֣�R���{����  0l�"
����o�/����MNo�����ګS!�����/Ɛ�vZ��CU����   ֱ�B\Z.�B�+�[   ���6������:��;`#���rjz*�s�K6����`�OU���    ���I��yo�'rw   '�l����������'Ϯ�q�ܳ�x� ַn/�>\���ʹ��   �oa1�B���   ��	� �|��uJ�އ�dj2�\YN�� `���z����?���   FW�����krw   CG���w�~��/��Ɂ������Z �C���~h�~��u��|�   `�--����:�
   �� X{˝�k��c��(.xY߱-��� `�i-��_��O=�[    8y���s~S��C��   7o���7���S�n8?wl3ӡ�{i9����ee5�|1-��G��q;   ���i�����2w  @nNpq��t{o��!!��SN��?t �Cz������n��R�    �����;����w  `�s�;��uv�.w�y�;`���8���8��������~t����V���    �B����l��   64'����^y{��(6��⊋��� ��jJ_z��=�h�:w    ä׋g�O��~���  ���~F�f�_��^��6�X�p�UE�,B�����1�o>�V���z�+��   ��������  ldNpQK��K�`���r�ԭ��* �W��O=8�>�t�n   `��V⎹���¿��  ��7~F������n7���6�͛Cy��q2w �)��~4��ۇ��q;    G����)�  �F�Q����Bu�yE����f�!�n`�<=���B���N~�   pLz+q�b���!��#w  ���m_�s�=��v�����$��br��X�� `������?�x�1n   �x-��_p�;  �9�`�t��u�`#ؼ9��������py�PZ�̃u��K)w    �[��v,lY}m���n  8��F����٧���rw���E�jL�b� ��r7՟~�^��w� w    ���X�b0p  6��!KK��n����ʉ���(@1����S��}�j�   p�u{q�m��_��  �d2po����n/����n˦X\~a���@~��P��ǫ�������r�    0�:���r7   �L� #bq����0�b�E3�s� �Uz���{��U��vj;    kk�Ϻ�m����  p����;����n7���F�E��ĩ[c#w ��ک��}U�s_�zU��v    N���î  ����`����`�m�	�����; �&=�h���G����T�   `c���ٯk�)�  ��`����yo�'��p~�e�����Y!�n��kw�{j{m�   @&˽�)�  ��`����u�s7��{������F� N����G���   @v�^<��˯��  ���ֱ��n�r�[�<w��f3W^\N�� ��ZZ
�?�̩�U�r�    @!��n���   k��`[^�#�u�����w�r�����s��[m��.[�dɒ%��Y@�@&;�L��qlƉC���Y^7���5�x�C����`l��c�6ް1�E���:��s����	p{����9U��_�yҥS�o�
�٥w;���`FdY�O<��tӤw�EW�   h��;��~py�  ��d��R��a�� ;?uL��۳��[��� ������n��w�S�Ip�   �FZY�>��  `-���`�_BtU���|�^wAg1u ��'���?�T�<�|��n   �WS�َ���a�  ��b��B�~nx�J?\����.�lذ�Y	`�M�1���jp����h�j;    �P��_�n   X+F[ -�����\o�5r�iYw׎l>u k������T�<�T�n   �#�R�s������   k���e������ K��V�N.����K$ �+��p,�uۤ?�:u    �� |*u  �Z0ph�lX_Wױ����E��6m
�� ��C+���w&��?��Ѵ   �[�g]�_���  `����ҍ�ԃ��o��iu�	�s��l!u k㩟����N�;x(T�[    ���l0ʮN]  ���Z����VU4��5��!���b��,u �k2��{���wW��
1u    �����M��q��   ����%�����+�콩;`Z�;;[8�Ĭ����u��8��7U+O>ǩ[    `��!�����  `5���x�	����0��;.���ِ��Ux�.�׭Uo0u�    X+˽���bqV�  ��b��_�J�;�ˮH���v6t:!K���(�X���N����.�i;    S��c�d��  S���~n��Q8)uL���g�mgd�; X�<���j���$u    ��C+���]Zْ�  `5������oS7�4�t���;��; Xq��uy�U81u    ��IU/���J�  ������(���;`]�/۰qc�� �ؔ�P��I��e�S�    @����/}5nL�  p��n��"uL��7e�y{�� ��_��T�<w LR�    @J�I8�ǏW��   8V� v���;{�|w��F�^�/fY�Rw p���ŷn��2��1    �+E��+��z-  �j� �\�OǺ6��U�s{6��l.u Gg4
��o���Xc��    �c8
'o}��oSw   w����s�K�����0m�!{���� ���?}{�{��8I�    MT�?��  �X�4ToP�]���vXe���ٰa�3@=�t~�U�(���    �
zE����/u  ��2�h����8{���%uL��O�:����Sw pd�:����w�Su��    �oy�2u  ��2ph�Q�w���0M�<�K/�,��� ڤ��׿3�=�t�n   ���������[Sw   w��Y�1�z��}g��6�wd�'���; 8|?}6���M���rp�    �H̖�U�+   ���;@�84����B��&sݐ]tngC� O����㱼�Ϊ?����    �he����K���   G���A��r\\����is�����{ � �o��*�}�*c��    �+ֱӭçSw   )C/�����qؘ����͡�gg>����VC��[��O�Q�    �˽첫�^؜�  �H�4�r/^����/�lȲ��� �սx0N�~S���K�J�    �b<��y8�/Sw   	w����s�?*����0Mvn�涜�ͥ� ��=�t~�U�(cL�    Ӧ7�._Z��!  @kx�����S7�4�tBv�y�b� ^U��ñ�㞪��m   �5Q���Cs��Sw   .w���/���/�;`�\tng��̳@CM&����U��a�    �v�^���   ������kB�Y���o
������ ��~?T߸��=�\��n   �Y0(:����oJ�  p8����o��;oN����v�,��@=�|��I��J�S�    ���u����+Sw   w�Ė_�\Wձ���ř�gݭ[��� ��,��b��;��hb�    �5�������oM�  �Z����g6���w��i��!����b� ~Y]�x���������v    H���ܡ��Rw   �w��F�������0-���-l�:�; ��q��}�����q��    f]�����R�O�  �j����`Z�/�삽��� ��A�o�R��;&�[    �F����0�D�  �Wc�����./�ٖ�0-.���0?���)^:&߸��-��:u    �/�"�H�  �Wc�HQt>����	�g������h��>�߼e�/�S�     ��W�;�f�|w�  �Wb���gn\��׏��i����,Y� Bx�Gqx�U���q;    4To�C�  �Wb�������1��j8cK��C�!    IDAT=��l.u��˲�p,��AU�:u    �jVz���|�/u  ��1pXg�}1����~3uL�,�择; f]�!�zw5���j��    xmu����*u  ��1pXgeY^5��0���-�)�� �e�I���m���O�q�    ���:���W���   ���`����R7�4�_�{;�; fYQ��7W���I�    ��L&q�ǏW��   �U� �诗T�-�;`\�7�0?�Y ������N�;���-    ���;W,-E��   ��M
�:*���`�)�����Sw ̪�=�߼e�/�S�     G�,�i��C�;   ~��;�:�̍+�p~�����ِe!K�0�{*��_U��    ����?��  �����C�kb4ȅcu��YgǙ�\��Y��㱼��U��%    �j���^�.u  �?3pX�^��ƕ~���0~��|їE �W��x�CUq�U��    Xm1��+SW   �3w�uPo>�/&�����nǙ�ܩ'g�� 3&�y_U<�H�    ��� ��/}5nL�  ��;��8ԋ���.�C���Ά� �$�o��<��8J�    ��I6����/Rw   �`������oe�=u��ޝ��M�B'u����o�^���8N�    ��~�0u  @� k�?.�1�vCv����v�u2����'��>'�[    ��Qa��ׯ�v�   w�5���x��ޔ����¼���0��[�U���v    �1e��D�   C1�5t����I�Sw@�-n����B��YP����w�ދC��    X�~�-K7�SSw   ���`-���n������B'Y��i����T��X�n    Ҩ�8�R����;  ��f��F������(;#u�������_A Xc+�X}��`��   `ƭ��R7   ���`������.9/���� k��r�|�U�(��   ��a��ϕ�I�  �.w�5���z����f���u�o��Rw L�/��7o��G�S�     �q�>��  �]� k`y�_��I�mv����]oX+����}[ݛL��   �_�d����m�;  ��d��ʖ�b�d�N�m�����r��� k��q��;�~Uٶ    �u���_��   f��;�*;���x8�'��6���;R7 L+�v    �p�������]	  ��Xe�0����f;���N>1�� �F��    ���/����  ��1pXEW]_�����;���<��殷��v    �H���  ��c����I���k+��wd�'l�:�; ��q;    p4��E�˽�;  ��b�	�J���|%�,u�U�	�}��� �Ƹ    8Zu�y�'Sw   ���`���)?6��M�;�����7��V�s/�    Ǧ_�w}�+q.u  0;�VI���8u�U����q�`5={ �o�ݸ    86�q8��g���  �� �����zE�'u�վ���¼����r;    ���A�#�  ��aH�
�U��b��ڨ��y�]oX-Ͻ�7�^��   ���/��}�wq�  `6��k�{���;������ϻ��*�e���   �U�A��d�
  `6���?��xSw@�uCv����v�U`�    ����KKq>u  0����J?�a�h�sw��s�G �Ջ��;w�    kg<����ORw   �Ϡ�|����EvN�h������'w��Z�շ����q;    ���E�"u  0��������C�����=�B��Y�X��b��۪�hh�    ��� ?����=�;  ��fTp���b>(:�H�m4?�}�\o8�"Tߺ����   �uRǘ�q���;  ��f�p�^��<�Sw@�N��v�cP���֭�~Q�:u    0[z���KK��<  ����(�'��n�6ZX��]�B����B����^�o�    ���(�|(�/u  0����gol[d��6:��B��� m4���[�M��V�q;    ��p�4u  0�����q�c;�;�m�B�w��� G��C���&���B��    �m���K7�SSw   ����(�E�ݩ���۝��pb�wU���I�    ���s/��?O�  L'w�#�7K廋�>=u��\7d{w��; �&�B��U�g�q;    ��Ax�  `:��ޤ�h�h�sw�ݮg�#u���|��8J�    ��e��oo�5u  0}�� ��5_���A����6�n����z;��z�X>�h��     x9E?��  �>� G��?6�����6�vw���=w �'�������     �de�}�W��Rw   ����E����6�N���Rw ��3�����_�N]    ��F����gF���   ���;�a��bg�����{vXذ���p\�[���    @��pE�  `���q���M8"�N���q��0�P�t{՟LBL�    p8V�ז���  ��0�8Le�����6����]o8<�Q��}{�/�h�    �F�C�P~"u  0=� ��ׯ�vQ֧��6�;!��6�� h���;߫��+�N�    p������  ��0p8������6go��[�<k ���ݻ���c�:    �h�쬿�B�M�;  ��`t����|��ޒ��$�C8Og!u@�y_U��8I�    p,����  �t0px/e�G'�p\�h�[���C'u@�=�x,{2�Rw     ��A�7��Z��  p��^CYf����<��^�O�������     �a4	��=\|0u  �~� �b��xj���O�mrƖ�{�	�����.�ɭwWE�S�     ���0�<u  �~� ������:��8����v�W1(b}��U��BL�    �����W-��9u  �n� ��濛����C��S3_
xU��߫�E��   ��3��|�o���  @����+o(v�lw�h��vbY��&�1�[��/
U�    ��2,��S7   �f��J�����N�a:~S�o;#�K��Tw�_?{6NRw     ��~�����Rw   �e�	�
�"\�������B����G�����(�Rw     �����ް�g�;  ��2pxW/�^W�:[Sw@[,nȲ�gf�; ������u��    `����S7   �e��2&u�㱮]���t�|!�]o�U�^�n���:u	    ��)F��}�wq�  ���^F~#u��\7d{v��� M3���;wV��(��-     �)�uV���  h'w�_���]6�SRw@[�ٕ�w�2��~Y��j���v;    0�V��  �v2p��I�é�-�<�}gw�Sw 4ͽ����$u    @*�Q8���л,u  �>� �����N���z�h�����7�N��&y��8|��j��     ���q1  �����mM¦�����,�n h���]�WE�    �&�ٯ_��X  pD�~���>���b˩�{�	����)�a�o�^5���%     �0��M��ޟ�  hw�����q�_�O�mq����Y�!�rg�/�P�n    h��đ1  ����\|��7�*nH�m���,?����v������8�bt�    �W��K���|�  �=�~n0�~ӹ��C���	{*�Q��     h��$.�F��  ��� ���/�R�Sw@�/�l��̕������"u    @�����n   ��� �0����c7u�����B'w���������J]    �l�~��/}5nL�  ���;@aeߓ�ڠ��]����̋1�[��2��-     M7����O�N�  ���;0�>��⬢����68k[�߰��྇��a��    �-�q���  @;�3�.�W���þ�;��3�g���Ï�a�    �6)z����ON�  4�A'0�E�۩�N;%tO���; R�����j��%     �Rձ��r�'�;  ��3pfڧ?_�+�|{�h���\of[U�x��&��$��-     m4翛�  h>w`���!�,u4�←oߚͥ� H�T��C�J�    �V�~v��K/���  h6w`��Exg�h��g��Y|�Y�=�O<G�;     ڬ�c7�,~$u  �l��̺��rOQ��Sw@��v��ϧ� H��J�.Rw     L�^Q�'u  �l��̊U������vn���=3 ���C����_U1u
    �T(��^z���  @s�3���L� m������̺�88���     Ӣ�c��?��  h.w`&}r��=(��;��N;%tO���; Rx��8�я�q�    �i3*�{R7   �e�̤n�>B�Rw@����z;0�������2u    �4���^z���  @3�3iXν3u4�←oߚͥ� XoU�w��Ub�    �iTձ;�H�  4��;0s>�T���Y�;������,��`��uU,��:u    �4+��  �f2pf�\�}4F�]x5Y��;��� ��ɟ��O�Q�    �iW�:^�����  @��3���H� M���l���s0SE�*Rw     ̂I���+Rw   �c�̔��0�V�����t���]ofM���j0���:    `V���n   ����)�:�H��>x�o���Oͺ�; ����c��    `���⥥��  �K�<��2��R7@ӝ�3[�1d�; �ˁ���G�a�    �Y3��C��;  �f1pf�u_�'e�7u4Y���]��� �e4�w��N]    0�&U�}�  �f1pfF1~��c7u4�Y������`6dY�w�WE��    �����ϧ  ���`f���ݩ���ٙϧn X/�=G?�i��     �e�I��}��  ���;0����"^����B��3�r ̄A�{���     �PT�S7   �a�̄'�,?TUa!u4�9gw\ofE���j0���:    �zE�ͩ  ��0pfBQ���n�&��l癙�;0|�x1V�;     �?F�pҧo�-u  ���Ի�k�S�ץ�&۹#��tB��`�\���?���     ��Q�_��  hw`��|p�{�qؘ��l�Y�ہ�c���[j��    g0�\p  B��('����N:!tN���; �ڽ����`�    �@�0��W.H�  �g�L�Aٽ4u4�n�ہ��a�ȏ�0u     ����^��  H���jW/�^W�)�;��:�,�ڞͥ� XKU�m�N�X�.    �����  ��܁�6�;����ma���< L�{�W�`��    �_�?��e�  `��Sm8�ޖ��l��|>u�Zz��0~�8J�    �k�u��G�W��   �2p����ckYdg�:~S�O;%�� X+�q���;)���     �1��R7   i�S�w(�H��9x{vv�cY���r�u1�v    ��⥥�W� `�~S��w�n����vn��� 0��{!��q��     ��L���`�7u  ���;0���r\,�����T����6,x ��d���VEt�    ��&���  f�a0�z�'Up�^��r����Cu1�v    ����S7   ��Si8�7u4��,;㴬��`-x1N{*�Rw     p�p�_�o�  3���J�~|}�h������,u�j����~=�n�    �^U�J�   �a�L���/�5��ͩ;���:3̧n X���*Wz��     �`4oM�   �a�L�b� u4�)'e���:�; Vۡ�X=�x��     `uE��ڥ�-�;  ��g�L�rޒ����r�ہi��~=���     ��:�|�����  ��3p��ҍ��r�J�M�wBر5�K���z<_<��    ��h.K�   �?w`�,�+j�m𲶝������ �K����e�     Vߠ�.^Z�>� ��M 0U�2�V�h��w�� V۝�UEU��     ���8l<��3u  ��܁�q��bgPf��&Zܐeg��uSw ���~G�<'�;     X;�x��S7   ������/�����D;���,Y���2�����u��    ����7�n   ֗�;05U����T���� Vӽ���(cL�    ��*˰��7���   ֏�;05�a���2N:!tN؜uRw ��^���G�;     X{1��W�J�  �w`*|��YE�oM�M�k�����1�;X�.    `��exG�  `��S!���b���&�C8k[>��`�<�X=\^U�     �OYf\��� `F�Sa8
oO� Mt�)YwÂ��P��z���0u     �k<����/K�  ��7����b^�y�;��vmw��w�_�Ub�     �_1	���  X�@�-g�oM�p\�h�N'�N�; Vó����q�     ���7�n   և�;�z�q����Dg��sY���X�����E�     ��qǵK+[Rw   k��h�b.M� M�s[>��`5<�X=\^�u�     ҩc�'U��;  ��g���g>�|JYf;Rw@��uC�uKf��^Q�z�#�0u     �u���  ��3pZ�?��@]�N�h���esy�� ���b2	1u     �����  ��3pZm<�����h綎��@�=�|���q��    �f�����oH�  �-w�Պ����+7���SB7u���1�{���     4L����	  ��2pZ�/�.�≩;�ivn��BY��c�����J�Sw     �,�q��  ��e��֠�|0u4��m��� �b4
���e�     ��(�=�^����  ��1pZk4oI� Ms����tB�� 8?�aU�F!��     �y�*΍���{�;  ��c���W��evN�h�gv�bY���uh9V�=G�;     h�:俕�  X;�@+=���eURw@����S7 �{��X��     �Ɋ2�>u  �v܁V*���n��9~S�OܜuRw ��<G�<'�;     h�r�o�vieK�  `m��T�R7@��8�3���h������     4_c>ʺ�K�  �w�u��ոq0�v�9kk�O� p��Q��B��    �v����  ��a���S��?��I�M���,?as��h��$��?RSw     ��(�(u  �6܁։1{g�h���f�����#�p41u     �Q���O�ܗ�  X}�@������4����R7 ���#O��    8b�(�7u  ��܁VYZ�[�avF�h������:�; ����ʪr�    �#7���n   V��;�*/u�c�Rw@��83�O� p4^:&O�4�Sw     �NE�]��  X}�@����7S7@�lߚͥn 8��N]    @[�&q�_����  ��2pZe8��>����g�	�g�� G����s�$u     ����n   V��;�W�P����Sw@�lߚ���Q��CU�:    ��+'���  ��2pZ�;���:K�M�����h�'�����P��     ��Eػ��_  `�x�Zc8�ޚ����B~򉡓��H��}W��     L�I�t�7�� )_�i    IDAT  V��;��a� u4��3���_5 Z�'��`��     L�Ѩ��  ��1pZ���=�Q89u4��3:�� Gb2�q��u��    ��RN⥩  ��c��B>�ߗ��d~!d��܁Vy��8CL�    �ta��R�� �)��h�a��%u4��3��B���p�F�~��z��    ��3��q�n���  ��0pZa8��O� M���|.u����h5O\o    `m�F�w�n   V��;�xW]_���ɩ;�):���~j�M�p��2֏�(��    ��)'���  ��0p/��K� M�팬��!K�p�z4�U�x;     kgP��KK�  ��{��uxk�h��g�s� WQ��ѧ�Q�     �ۤ
��śSw   ���h��0?7u4E���uK�M�p��?R�u��    �Y0v~'u  p�܁F�ji�}4�ON�Mq�)Y����7��"֏�8��    ��(���  �cg 4Z����:K�Mq���\�������     ��a��K�   ;w���exk�h�3�Ȼ� G����    ��F���?�����  ��1pm8�n���||�o\�� ��V�X��     `�,/W�N�   w���^z���0?=u4Ŷ3�\���1(B���]o    `��F�7�n   ���;�X��q�c�:?w���h�����    @�q</u  plG�����n���_٩'g�� ��(c����     $R��S>{�`[�  ����5f�n��8sK�B�Rw ���e]��     `Vź�V��ݩ;  ��g�4��oqa8�w�8sK�K� �Z�a�{�v�    ���Ix[�  ��c�^v,;���ڻ��]}��A���%� ;��8N��A�K�E�� �� ����2�P���(���A)�M6�fX]{�/�PdQ���~���y��7��U]�_�8w`���_��ˡ�etLAnRz�n������Ѱ��    �̭V�7�  ��3p&�,�(���\.=��i[���͛��v     �����ע;  ��1�&���w�`*^��w� ~��~���!9�    @��R���qt  p1��$�����0��m�� �L�������    ���5�4�  �w`r��ɳ�u�0���� 5GGi������j[��    �����ft  p1��-�(� ��{��v`�jM���z;     �r��_99�v1  ��� LΪ/ߍn��x�N�� �˼�Nm����     ��~HW>�;���  ��܁�Y��_�n�)�MJwo&܁)��ò��     ���t��   ���;0)������k�Fw�ܹ��˝��; ~��j��iu�    �I:[�ߋn   �����>��q���&H)�|o�z;0i����    0]m���  ���H�Ii���`*^��v� ~����:Dw     �/rv��~��7� ��1p&嬭�� S�%�ײ�40Y����v     &��U��*�  8�9`2NNj�j�ע;`
^��vjM9���<}V��>�}t     �*5-?�  8w`2��N���u?����;�2�����U-�     ��"  �����[�atLAnR�w;��Զ���Nj�;     ��x�j^;9��1  �A� L���ntL���y���L�~R�a��     ��C�;�;�nt  ����Ѷ��0/�i\o&��T�f]Ew     �y����� �1p&�7�������{��Nt��y�~m��U��    �(C�;�  ��܁I�GGXK]Dw@��"��׳����_�ph�;     ������  ��3p&��?�n�)�s+-�&���������$�     p^������;  �/�����[�ftL�Kw�et����7�*�     .���X^��Ϣ;  �/�����6}-�����l�L���4��A�;     �κ��  �!܁po�<��j��������㴈� ���歡�%�     .���   |1�@�U��*���; �K�]o�o��RR��۵��     ��j��F7   _��;.��?�n�)�w�YF7 �}oݯm�J5�     ^D�77ON���  �W3p����0{�`R~���z;     �����  �j�@��˯E7@�����Et��k��q�;     �2�����  �_���''g_k�z��^��z;0=�VYE7     �e����  �W3pB�7�_D7�ܻ���r�J����     ��r�j�]  6��;j��ߍn�)�}3����;�-Ct     \��-�����K�  �/g�����p��գ��_ɞ��d��<��     p�J���  ��3�B�V���g���r�����٧�Dw     ��[z�8  L��;�_���_m�z����j܁I������     l�UW�e  &���̋� Sp����t��R��~�;     `m��Jt  ���a���^tD;:L��~�<&�Go����
     G��k''�^��   ~1�: �j����ٻ{;��LI��K     c���O��� ���a�6�� ���4p��jz��o    `�u]��  �_���'�_j�t����n� �ͷ]o    `�u�x�8  L��;b��� �R�%��ж���v�     0���Jt  ���!�.�ntD�w;/� ��[�     0�U�o��y��  |>w D?ߌn�hwn5�����;��n     �������?��   >��;b�.�� ���p���G�S��qr�    ������� �D�k��'��.y������ё�00o�]]o    `VV%};�  �|�u��.��I�)Gw@�;7�ҿ`
JI���C�     ��u���  ���k�|��atD�}�YD7 �����k�T�;     `�V]s�{߯>� �	2p֮�oE7@�;7�2� ��~�vi�     `��Pw^}��w�;  ��g��]�*_�n�H�"����5 ��*��?�}t     DhV�ߏn   ~��;�V''�i��RtD�u=-�&����߭m-�     �m�oE7   ?��X�g;�o�Cڍ�H�o��LÛo]t     DY����  ��3p֪+�+ޘ��7�et��'ux�8�     �[�/E7   ?��X���^���ݺ�;����n     �Hm����<}5�  �Y��Zu]��7f��Qn�v=�X9���wk�     �>���  ��e`�U�6�D7@��7�2�����?=M%�     �u�ߌN   ~��;�6���ö�7�; ���"�������     �R:үE7   ?��X���<�'����n]s��Uk��[�     ��w��  �g����D'@��"�k�ٳ������T�;     `
�nq���  &���ڴm�vtD�u#-R� �O�-��    ��ꇲ�����  ���;�6�!�� �n�ȋ�`ކ!��j�     S��y���  ��2p֦o�������������T�;     `J��~'�  �)w`-�8yz�����t�ZZF7 ���wK�      SS����  �܁�����RrtDٿ���~����}*�}P�    ��i����  �퀵(��NtD�y��v ���+Ct     LO�6w������   >c��EߧoD7@��׳_��~�nq�     >�P��տ��  |��X��K�E7@�[�@�����G���     ���y�nt  �w`-�>ߋn�(�I��5w ��RW��
     ����ߎn   >c������t�Q�r����y��E7     ���Cz=�  ���0��;+�rc�n�h\o�%��>�}t     LY��W�  ����;[�ߊn�H7��et0_�_�aH5�     ����퓓jG  �s`tCm�� �n\�.�a�yP��     ��~H�OvW>� �	0pF���+�%7)]?Ξ�@�ZS}�A�;     `Ԛ�At  `�����/E7@����,���@�־�S��     �MPW�ף   w`d��u���qtD�y=/���z�A�     `S�����  �������+��^�l]���!rN�����;     |A]���   �#r�����q2pB<|T��g�Fw     ����|7�  0pF�v�[���q6pB�w�     Υ����ɳ��;  `�܁Q�}~-���fo׳��΃��n     �M�,��F7  ����j��JtD�y��v ���4<y���     �4mͿ�   sg���7� ʍ��@�����     peH_�n  ��3pF�''g_뇲�Qn�1�_��     �Dm���   sg��f/�� ��'w`��>�V�    ��.ߋn  ��3pFS��[�ew/��+�sX�־��
     �L���:9�>� �@~ F3��k���qv��އ��v     ��2ԝ���W�;  `�܁ѴC�jtD�~�܁��9��ޯ�     �)�Nt  ̙�;0��o�E7@�kǍg,�v����Y*�     ���P��   sf|��{߯��M7�; ����w`�|�z;     ��a�_�n  �93pF���7K�����������;�v�?�    ���jt  ̙�;0�OO�w� ��An���;�y��T>z��    ��}})�  ���EߕoG7@��Ǯ�������]     ���7����3?  b��b��W� ʵ��]�ڽ�aq�     .A-u�<�Vt  ̕�;0��4^��l]��=_��{�a5p    �Kr�d���  0Wx�(�>݉n�(ׯ���׳gi8=M%�     ����  0W��(���� ��=_��z���     p��:��   se�\����/u7�"\��)�����w     �DmM�D7  �\���J)�� Q��Et0;���.�    �e*��nt  ̕�;p�ڔ�� Q��6���Z}�I�6��     �&m�nF7  �\��������r��w`�����v     �l}_�O�k��  sd�\�a��D7@�����
�Ճ��;     ����ߊn  �92�.]��{��Y�tx��
��PR��Q2p    �t)�Zt  ̑p��6yM�tt�)�����G�/Ct     l���_�n  �92p.�o<8l�|��_͞��Z}�Q5o    ���R^�n  �92�.�����H��`�,�Et0/|\��     �V}�_�n  �92p.ժk~-�����Q)�>|��    `$}�oE7  ������ztD�z�\p����C��     ���������  ���!�T}��� r���#܁���a�     `��R�.Ͼ�  sc�\��ԗ� ��~jM���||���     ������  �w�R}�� �]u�X�ZS}�(�    ��V)}-�  ���TÐoD7@��Gi� ���Gu��     [o����  07���99��]��; ����3X��%��    `��jt  ̍1pi�����V�W������>�6}\�    `�>ߍn  ��1�.��Y�ftD9<���`rN��Gu��     �9�K��   sc�\���ף �b���~���<<}�J�J5�     �����  �w��tC�rtD8<�����;�?�}t     ��0����ZoGw  ����������0{�k���e�n     �9yr����  0'y��)]�W���ѡ�)�>}�\p    �5*i���  ��<�ҴC�� �6���Z�]*O>�%�     ��×�  `N�K3�jtDp�X��?��y;     �W_�K�  0'y���w��ɭ~H���� -��yx�q�     `n���E7  ����b(˯G7@��"�����;�y��q�     `nj�oE7  �����ˋף ��a]��܁����O\p    �uk�t#�  ����C7�� ��g)�����Z��     s3�Qt  ̉Qp9J�JtD8<�,���#��     B?�����܊�  ��0�.E;����p�w`=>~\�     �P�_�n  ��0�.E��,���;     ������  ��<�R�C�� �x��5Տ?I�     ����  ��<�R�C=�n��������<�eR��     �����Jt  ̅Q������{}���;`�vwS^���l�O��>�     欯�nt  ̅�;��~���~5�j���d�Q`->~\Jt     �Y���  ��<�����E7@���Q`==�Ct     ��P���  ��<��������`��CΩ>z��     �04G�  0�y��5�3K����(0�g���}��     0g��ON�� `����~�w� ���:<����     �J������  ��<��eq+�"�{��{�$�    ��O���  0�y���܈n�G�sݣ���     &�-���  0�y�Js=��mw/��"��`�}��w     ���^�N  �90p^X�ի��n�W<C���T����     �4�^t  ́q�BNNjӕt��v��]oF����     05݉N  �90p^H{��^-i�붿�
����R�     ���C��   s`����i~=�"�_ɞ���?�.�    �T�zt  ́q�B��^�n��Wr�n ��'O��;     LDW�qt  ́�;�B�!�� �\�ƕs�����     |���at  ́q�Beq+�"�#���֮O5�     ��P����_�  ���ҥ���Y������i�     ���5�o��so9 ���/d���X��e�˝��;������;     LM�ҫ�  ��܁RKs-���`߸ߓ��D7      ?���+�  ��܁2�t5�������S�    `rꢹ�   ��@x!Co���\�����Yu�     �fH��  `��/��|� �����v[���m��     ���|3�  ���;pa���ם~�W�;`ݮ������     0I5Uw  ��pa����Z�K��Ε]_����|���     ��u�^�n  �mg�\�N[_�n��.�#{����     ���8�  ���pa}^�� �������>s�     ����Qt  l;w��j*�� ]�O`\O�U�    `���F7  ��3�.nHw�`�����;0�ZS}v��    `��R��  `��VJ�� �v�o����4��    `�jI�?=yx�  �����Z�k��nW�<;�q=;5o    �)��=|)�  ���pa�.�F7��]��.��z�i2p    �	[��Nt  l3w��J��������էϋ�;     LX���  Fd�\�����X�ݽ��	��w     ���mnG7  �63�.l����ٹ��]pF���j�     VR��   �����24���nWv=;����.�    ���1p ��6���ٹ��\pF��,�aH5�     �%J=�N  �mf�\ȟ�y�J݉�u�]fw`4��V��    `��� �����    IDAT�܁9{�z9�"�����i2p    ��+e��   �������r7��-7)����9}�;     L].�Qt  l3w�B�PoE7���|6n7pFszf�     S�׼�   �����!7ע`ݮ�f�v`T����     &��t%�  ���;p!C�7�`�vw\o���y��     �/Wjڋn  �mf�\H��jt��ޞ�&0.�    `����  �d�\H_�qt��ޮ��x�.��O.�    �ĕR���u?�  ���;pA�(� �mw�����j�     ���Vt  l+w�B�`�����5��h����      |1{;���  ��܁ɹ9�n�us���;     l�����  `[�Rj>�n�u�3pF��y��     �S�ō�  �V����>�3;{����x����     �!�"G7  ��2�.��u?��m�t���d�     ��V� `$�������`��v�ہ�<?�5�     �b����   �����Zܙ���w`<g��;     l�!Uw  ��;p!eH���n;Kw`��zֺ�     �I�	  ��܁s;9��P�Nt��b�r���8�V�V��    `c��� �H܁s{�>>��Зy���5��l���    `�)�G7  ��2pέ�rp=��mwǾ�٪��     �J��   ���8��Es� ��;0��6��     d�u/�  ���;pn���Zt���;0�U�\p    �R��  0w��J�� �k��h�*�     �Ajɻ�  ��܁s[��8��mgi���w     �,�Խ�  �V����|� ��;0��*��     ���5�D7  ��2p�-��jt���2��9[��     �����   ���8�E>�N�u�Y���笭�     �A��\p ����6�t� �Xڷ�Y��     ���89q�  �`��[S��;��l\p�1�T���     6ͳ��zt  l#w��jJ�
��Y,܁q�m5n    �t�XF7  �62pέԺ� �\F ۪m]o    �Mtu�ߏn  �md�������w`$]o�     ��v��  0w���`���4��;0w     �Lg�b�  #0pέ�l�����ط�h;w     �D;)_�n  �md��_u���Y����m��;     l��4.� �܁s+��D7��-�����    `�݅�  0w�ܚ�ܙ���w`]�;     l�UُN  �md���P]pg^r�R���8V��     ���"��  #0pέ�d�ά,�v`<}o�     �(7��  F`��[M�2��i�4p��u�     ��j�;  ���8�R����ҟt #�w     �D}S��  `��kZD7�:5�w`<�`�     �(���   ���8�����i�j����]p    �M���]�  0w��j���Yi�v`<��;     l�a؉N  �md�
�_���yY,\p�����     6�r�s  ���s+�w03M�oFS���     6Q��  0#U��\pgf_��H�!�      ��Z�2�  ���p.''�)�����4Mr�E�'��    `C�\� `F�������+֘܁��b�     �*��"�  ���p.��O�� �X���c��    `S��;  ���8����^t�[c��d(�     �E�Z� `�����b7��m�x\�(%9�     �ִ�n  �md��Ϣq���i�w`�w     �X9/� `���\;�.�3;ټI�.�    �ƪe�   ���8�n��:����%0�a�.      .���;  ��b8�ՙ��3?���HJq�     6�_� �8܁�9pʚ���E)�     �E55�  F`�
�K���3?�ꁑ��     l0�$ �܁s�2�Et��� cj�p    �U�7A �L����}���[)`4��     ���� `������?��Oξ�qط    ��A"  ���8���s��R�Hj�.      .���O `����4��@g~|��q�     6U��� `�����~� ���0�j�     �f�  `���,���O��/��Q�    ��9"  ���8�R�"����`,5ew     �P9{4  ���8�!: ����u;     l�Z�O `����f�?�       ���� `�  �	w        ��           L��;           �`�          �$�          0	�           L��;           �`�          �$�          0	�           L��;           �`�          �$�          0	�           L��;           �`�          �$�          0	�           L��;           �`�          �$�          0	�           L��;           �`�          �$�        ���{[n�:�0���h��%QQ,˒�����'N��Ԉ�H �F�b*)�#;�Lqok=�����{ @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @�           DA�          @��       w�K�z7�~M��4�7�w    q�     �AH���"/��<�������tz�
�   �[z       p7��7W�`V��    �K�      #�N�/�lX�^    �C�      $I�6_�=O��	�    >��      L�����^/�Bo   �O!p     �4�O����e�    �)�      p�F�G���lz    |,�;      �����p�xz    |�;      �y��u6��w    ��#p     ���t'�7Y6.C/   ��"p     �#�$i;_��H��	�    ~��      �D�����y��v��    ���     �����r���2�    ��;      ����v<{~z    ���      ��tz���C�    ���     ����/��|z    ���      ��|��2��e�    ��	�     �%I��ޞ�i�	�    �      p�Ҥ����{���   ��&p      z����/���   ��&p      z�^�7.v�����;    8^w      ���ӳ�h�xz    �I�      ��Y��j0�w�w    p|�      ������Ȳqz    �E�      |@��oΓ$kB/   �x�     �J�As��O�$kCo   �8�     �_�e�jv��2�    ���      �M��b7���
�   ��'p      �����z4~�
�   ��&p      >�,���`�oC�    �p	�     ���/^_f��>�    ��      �I����H�~z	    �G�      |�4�7'�o�%Iֆ�   �a�      �,�&����e�    �;      �Y���n���}�    �;      ����'���U�    �;      ���?^��6�    >�;      ��ח�`��   ��M�      ܁��o��tP�^   ���=   �w�d�ywҶUz	   �e:��M����;x8�$k�ӷ���w]�-    >��  "�4����OO����  �q���p-n�sd٨����X�������{    xX��   ��nߝ�\}�q;   �m<=[N��V�w�p�y1�_\��   ���w  �L�V�z��'M���  �������7�w����Onۺ���E�-    <w  �Ⱦ��nW��U�5n[  ��ǧ����S��3���eӖ�j3�   ��A4  �&]���ds��Sq;   !��v��zz�'?y�>�O��w    �0g   ��\�o��ㅓ�   �?����e����Oߞ�ٰ
�   ��	�  ��K��?]����m�,�   �S֟�ONߞ�zIz�+M�6_��H���   ��	�  ���ӛ�O����"�   �W��\��=ɲQ5?yu��   �o� �=��7���e�4U?�   �W��Gz�:Q�{4��4qz    ��  �}��d�]N���  @PI�5'�߽K�~z�g<~r�6e�غ�   ��OX  ����A�[M��MBo  �%I��oγlX�����^,���W��Y�-    �%=   Z�&��r��.��v   �K����y�?-C/�����l0+B�     .w  �B����^�uUBo  �^/��o/���>��?Iw�x}�f�*�    �!p �/`_�ǻ�լk��  @f������.���$��|��<I�6�    � p �;Եu��}?/��Q�-   �����G�G��;�C�lX�ߞ�zIz    �	� ��������2o�*�   �a<{~=?��~�`0��//C�     <�;  �^]�l7W��X�CO  ��O��L�g��;�c������ӛ�;    �z   <duU��j�umz   ��h�x=��X���b:{�l�*+��<�    �� ����d�[M���   �4-6���U��9��7W������my    G(=   ��.������  ��.?y�>��|I7_��H�az	    �O�  �`_�ǻ�լk�$�   ��l0���^�zIz�i�����y�dM�-    �/�;  |��m����y�ߌBo  �ɲq�/ޜ�z�����e�:?}�    GF�  ��~�ݮ/򶩲�[   �C�lX�ޞ�Iֆ�w�ߟ�g����w    p�  �k�6�n�fe���   �&M�M�x{�&�&��F�G���lz    ��z   Ĩ��A�[M��MBo  �_�$Y��~�.ˆu�-�%Mg�o�����Uz    _��  ~�k��n5��bz
   ��$I���ͻ,U���}��__7�~PW��   �4�   �E]�����\�  @��n~��E�?-C/���t���E���   ��	� �����x���um���   �-��W�a^�^�-I�6_�=O��	�   �/C� �Q��&�ܾ����(�   �������bz��e�:?}s��%]�-    �=�;  Gk�ߌn�y�TY�-   �1Ƴ�����M�Z�?-g�o.C�    ��	� 8>]�l7W��X�CO  ��5��-�ӳU����t;��-C�    �n	� 8*uUnחyS���[   �c�Ə�����; 6���l0+B�    ��5���    IDAT�z  8]��v�I]��S   �Sǧ����U�����5��-}    D� ����_�Ӯm��[   �S��v��zz�h_�L��=	�   ��%p �����oF�w   ���fE�x}zĨ*����_���   ��� p���I���m�,�   �TY�?9}{��%]�-��ތnW}��un�   8@w  �~���zz   |�,���>�i�����g]פ��    �e� 8]ۤ��ͤ�KϹ   <Hi:��Go��$kCo��4M�_]&n   8l�  B]�b��t]�jj   �4�7��w�Ҥ߄��i�*[/8�&�   �/K� ��ֵ�n���U1=   >W�dm~�ݻ,֡�@lڮIW��ڶ�m   �x	 ��U�e��.�Nm  �aK�����,U��@l��M��?��M�p   �#!p �A��q�ߌB�   ��'��W��|z	ħKV7~�4�0�    �� ��k�t�]Nۦ�Bo  ��k���r8\�B��t�z��ӦڌC/   �~	� x0��ͨ,�>j  p����G��m����_����$�    �� ��um��v7��.=�  p&�����W��w@�n�{\�7��;    C  @���դ��$�   ���ӛ��lz�h{��Ӳ��C�     �;  q��d�[M���   we4~���^,C�m7��(v��;    K� @t����ԩ�   ��h���/�B���y�}wz    �	� �ʾX���fz   ܥ� ��'�^��1ڗ������
�   �8� �B�V�n���M���   w)̊���E���\�77{z    �� �~���zz   ܵ�?ٟ,^_�zIzĦ�nG뛿<���$�    �!p  ��m���f�ԥ�R   N�����E�dm�-���oo���k��    �!  A�U1(v�I���	  ��I��99��]����[ 6MS���??�&�   ��� �_]��v�I]��S   �KH��=y��wi:��/�m����?�&�   �8	� �7u]���r��v   U�dm~��]����[ 6mWg��g][��   �Uw  �žX���fz   |9I7_|{��O��K 6mפ���|�6�[�    �Mw  ������v5i���\   ���/^]�}�%�.Y/��Y���K    ��� �/f�ߌ�b=�   ������p�؅�����ǧM�s�    E� ����&��n&M]z�  ��M�/�F�G��; F��T�zz    �� �;UWŠح&]�&��   ��6�=�O��C�ݮ��*���;    xX�  ܍�Mv�դ��A�)   p�ӧ7���*���f�ߏ��zz    �� �߭��~�]N��  ����Ng/��w@������˓�;    x��  �.�b=.��Q�   p_�|;ϿyzĨ�^���bz    �� ��ҶU�ۮ&mSe��   �}�fE�x}zĨ(�f�����   ��&p �����QY�ǡw   �}������^/�Bo�����t��ۓ�;    x��  |��m���f�ԥ�H   �J��˓ś�^/��/T�z���I�   ��& �Q��դ��$�   �Oi6��Goϓ$kCo����f���˳^���   �;!p �um�ۮ&u]BO  ���$Y�/ޞ�I�	�bS���z��^ρ    ��;  ����~�]N��  �1J��=y��wY6�Co��4M�_/����4�    �� ���q�ߌB�   ��$m��7�lT���i�:[/8�&�   ��#p �_�m��I�T>P  p��n~��E�?-C/�ش]����?k��wF    �/�  ���~3*��8�   i�xy9�E���k���gmSBo��e�N��6u�g
$e[�w:ޞ��Aql'�x�[$!� A ��Nw:���]Ej�+x���  p�� h5u��l�j��}  ��6ʾ~�Cw@|�d�x}^UE/t	    �̀	 ��ۗE��,�MS'�[    �����`��.tħI��볪\�C�    p�� N6��p�/�R  �{o0���F���|��QY�Cw    p?� �C���S��#��  @��<�G�ǋ�������n9
�   ��a� p�l�|�ۮ�N   Z�V�?]��'Bw@�V�O��b~�   ���� ����2ݬ�ú*��-   �n7�d�g7�; F��Ͷ��$t    ���; �=�ۮ��"��   �Xt��"�=��1*6�Y�����    �~2p 8bM]�7�Ű��|�  ��H;�m6}~�j%M��MQ|���=�   ��e� p��e�-6�a��I�   �E;헓�˫$I��-��n>Z�?>
�   ��f� pl�:٬�����N  ��$�N59��Ҹ�U������    g� pD��]���GM��v   �GI�V��7��S�n�ؔ�]?_�9o�gJ    g� p$��rX�ֽ�   �$I�l��*M�e���~���-��   w �W�e�^�GM]�C�   @|��d����B�@l�j���ϛƹ    �0p 8`��-�A�   �SҜL�^w�'��%��.����E�Ti�    �G�  ����f�V���9   �7�ٓ�^o�	�������w�ԥ�%    ���
 ���ˢ[l�æ���-   �Q������:tĦi�v~�ꢮ���-    �K� ES'��r��.  �WǏo�Gw�; >M�\�>����    �w ����:�f>jj��  �������2tħI�����\�C�    ��1p �\�Y��ګZ   ����h��<t�(_�}T��0t    �w �H�u��W�QSW��-   �n�gO>�������(t    ��  �mW�m�Bw   �!H��"�<}�b����t[ܞ��    ����  "M]�������4t   ��3�Ng/�Z��	��Y��>�nn&�;    ��0p �ľ,��f9l�:	�   � M����U��6n��)6�Y�����    �?��  ��N6��p�/��S   �P��^����J����)���ݻ�;    �c� ���:�f>jj��  ���nw�l��t��-��n>Z�?>
�    ��  �b���u/t   �$I�l��2M{��-�r��?�   p�� ���.��j>j��   I���ً�4��[ 6�~��o�[�Ɵ   8h�  _�n��o�|�   OҜL�]w;�]���~���͍�   8�  _@SW��z>��2�   �'iN�O����]���]'��>o   �8� |f���n��Q�   8T����t�bS7�4���h�ʣ
    w �ϥ���z9��n�   8T�����Bw@l�j/o�����}    GŁ �g���:�f>j�:	�   �j0��G�����������yX   ��c� ����ܭ{�;   �������"tħI���gUU8   �(� |"U]���|��U;t   ��`v7Ξ|��i�|��*W��%    �� |��-r�   �'u{��${�>t�(_~��,�a�    ��� �������|TWe�   ]����M���]��r���    ���� �#�ˢ�Y�G�;   ����v:{y�j%M������]�!�    _��; ����f���E7t
   �v�+3�v�E��ߧ���$t    |)�  �~���Ũ��$t   �v���������u��M��Ί��,t    |I�  �S�Y�ݺ�   �E�ݩ��7��S�n��Ň�z��A�    ��� ~CU��f55u��   �"I��d��*M{��-��n1\�?>
�    !� ���v��� t   ���fϯ:��.t	Ħ�������    ��; �/hꪽ^�GuU��[   �$����u�3ކ.����������V�IB�    @(�  ?�/��f=��   �c4�>���������v����ڡ[     $w �����f���E7t
   �Q���~�t�bSU�N>ua�    �  �V���﷝b�5u���   �Əo��w�; 6u]����E]���-    w ��ۗEw���Bw   �������2tĦi��r�ꢮKwv    �?�� ���گ�  �s���W�����w^W�n�    ��1     �Yt���8{�!tħI��7g�~�]    �1p     >�n7�d���Cw@|�$��9��� t	    ���     ����h�͞_�ZI�b�/�X��0t    ���     �d�t�˦/����_��N��b�    bf�     |�Wf�/��IZ�n�جW�f��f�    bg�     �i�v�ʦ/��I�
��٬�&��z�    ��;     �$IZg�o.Ӵ���)��'�����    �Ca�     |�$i����e����-��n>Z�{�    ��;     ��d����B�@l�]>X-~x�    ��;     ���d���ˊ�%����狷�V��n   �Cc�     �a������d�b�߯{w���Vm�    ��     �CF'_}�Bw@l�j���ϛ�r    ��     �F���,����}����i�4t    2w     �w�-G�ǋ���٧��o/�zo�    ��;     �z���8��m��M�T������uC�    �10p     ~U�7Y�dO߇��4I>��^�    8�     ���鎋l��&tħI����j��.   �cb�     ���;�Nf/�Z��	���o�e>�    ���     �i:�e��������|�    ���;     �O���>;}y�N�:t�f��t�+nOBw    ��2p     �O��U6�沝t��-����l[�LBw    �13p     Z�V��$i=9��e����[ 6��:+����    p��    �V��nN�ϮҴ_�.��Ň�z��A�    ��    ��K�l���=ن.��lw��u���    p_�    �=7���M���; 6�.���    �%�    �=6���ߛ�Cw@l��U?_�=o��$t    �'�     pO��q;<�����׽|��ժ��   �3p    �{h0��G������u����ܣ   @ �     ������E��M���|��i�4t    �W�     p�t���8{�!tĦn����ۋ�.;�[    �>3p    �{���6���M��M�T����E]�[    �3p    �{ 펋l��:tħI����UU�B�     �     p���p;�>�n��&tĥI�����\�C�     ���     �X;����u��u��M�x��,�a�    ��3p    �#�$i5�}s�N:U���]���r���     ���;     �$I���_/��q;��*��tW�OBw     ���     �L��u6{q���2t�f���ٶ����     ~��;     ��9�>��tF��%�b}��i�    ��3p    ���4'ӧ����6t	Ħ(>�׫wBw     ���     ��x��כnBw@l���h���(t    ���    ��N���Cw@l�]>X-~0n   �a�     n0~|;��; 6ey��o�[�&	�    �>�     p����ht�����׽��[�v    80�     p�z�ӻ���y��MU�:���y�T��    ��8�    ���e��?߇���u�.�.��JC�     ��;     ��;.����������wM]vB�     ��     H�m��W�V҄n��4M��o_]�ն�    �x�     p �t��L_\�Zm�v�'M�\�>����    �s�    � ��^����J���qi�|���*W��%    ��g�     �K��ʦ/��I�
���o���0t    �i�    @Ē$�'�//Ӵ���Y�?<,w�Q�    ��1p    �H%I��f/.�tX�n�ج�N���I�    ��2p    �(%����u�3څ.�جW�5�7��    ��g�     O���ˊ��bs��Y�    ��0p    �Ȍ����{�u��MQ|���=�    |>�     �����`��.t�f�[����Bw     ���;     Db0���F���r�V���Bw     ���;     D�?x��Ə�; 6�~��o�[�&	�    |~�     X�?]��'Bw@l��u�nn�    ���;     ��e�l��&tĦ�v�|���i*�Y    p�8    �@:�q�M������>��.��JC�     _��;     �v��l����J��-������o/��n    �<w     ���i���^^%IZ�n��4M��o_]�ծ�    ��     �����Of//����d�x}VUE/t	    ��;     |!I�V��7��v�
�qi�|��*W��%    @X�     �$IZg�Wi�ۇn������e>�    �g�     �]ҜL�]u:�]���*��A�]�Cw     q0p    ��*iN�Ϯ�ݓm������m�!�    ���     >����M�7ل�جW�n77��    @\�    �3ey�Cw@l��uV�/g�;    ���    �g0?�݅��Ň���݃�    @��    ������2t�f�[�����     �e�     �P� �����ؔ�|p�����j��-    @��    �����q��C���~���-��   ��f�     �@�;.�����; 6U����7�MS��    ~��D     ����p;���j��&tĤ�v�|��¸    ��:�     ����`7���j������L��WM�OC�     ��k     ��i��N_^%IZ�n��4M�^ο�h��cK    �b�     ���T���U;�T�[ &�3n?��m7t    px�    �J���f/.Ӵ��qi�|���o��K    ��d�     @���ً�4��[ 6���}���     ��;     �nIs2yv��v�K 6w����r�    8l�     �$����u���K 6��o��b~�    8|�     �;�&_����������l[����     ���;     �������`�b�^_N���4t    p<�    �WF���b�bS7'��李;    ��b�     �F� �/Bw@l���h���0t    p|�    ����q��C��M�����Bw     ���     ~����'����; 6ey��o�[�&	�    'w     �iw\d��7�; 6���w�x{�j���    �gc�     �#����˫V+iB�@L�j���ϛ�r�    |V!    ��j��^��ÿ��}����i�4t    p��    �����~r���v�֡[ &u�O���^4�޸    �"�    ����N�;�l'�*tĤi�v~��y]�[    ����    �{+I��d��*M{��-�&Y.^�WU�]    �/�     �SI�͞_u:�]��K���7gU��.    �w     9�>��t���%�|��QY���    ����H    IDATd�    ��3�>������������.��     �/w     �Q���~�t�b��:��'�;    ����    �{c8~|;<���Y��Ͷ��$t    ��;     ��`t��.��; 6��:+����     ���;     �@� ������Ň�z��A�    ��e�    �Q����q��C���vw;Z�?>
�    ���    8Z�n��&�nBw@l�]>X-��   ���    p����fϯCw@l��U?_�=o��$t    ���    pt�t�˦ϯ[��	�1��׽|��ժ��   �(�    pT�i��N_^����1��]'��>o���    -�     �$I�l��t��-��.�|��i�4t    ��1p    �($IZON�z���}��I�T����E]���-     ���    ���$i��^\�i��1i���߾���]7t    ��a�    ��K��鳫Ng�]qi����yU��%     ���;     ,iN�Ϯ�ݓm��K���7gU��.    �#�    8X������d�b�/�>*�|�    ��2p    � �N��0<X�����?<,w�Q�    ��a�    ���.��Y�b��:��'�;     >��;     �?x��/Bw@l֫w�mq3	�    �g�    p0z���8��m��M��Ί��4t    ��e�    �A��&��������0^��=�    �)�    �Nw\d�g7�; 6��|��|�    �S1p     jiw���^^�ZI�bR���j�q;    pT�    �V�v��q;�LY���ś�V�IB�     |J�     D����ӗW�$�C�@L��u�n�ָ    8J�     D'I�*�}s�N:U��IU�:���y�T�x    ����    ��$IZON�z���}��I]��r��i�4t    ��b�    @4�$��ً�4헡[ &uS����.���n    ���    �DҜL�^w:�]��I������E]m��[     >7w     �0�>����"tĥI���gUU�B�     |	�     7����;]�4I>}V��A�    �/��    ������݅��䋷���n�    �K2p     ���|>�/Cw@lV���r�    �K3p     ���A>��"t�f��t�-nOBw     �`�    ���OW��ɇ������mq3	�    ��;     _T��m�ɳ���b}���Y�    ���    �b���fϯCw@l���x�z� t    @h�     |ig��L�_�ZI�b��-����G�;     b`�    �g�N{e6{q�$i�bR���j��Y�    �X�    �Y%IZMf�\��N�b�߯����y��$�[     ba�    �g�$i59��e��5n�PU�n>7n    �9w     >�$I�l��*M�e��IU�:��o/��rO    �3N    ���d����B�@L�f���WMS��[     bd�    �'�4'ӧ����6t	Ĥn����ۋ�.;�[     be�    �'5�>��������������uC�     ���    �Of���}�w��qi����YU��%     �3p    ������Bw@\�$��9��� t	    �!0p    �O�����2t�&_~��,�a�    �Ca�    ���<�G��; 6����v1�    pH�    �h�^�>ɞ|��Y��t�->d�;     ��;     %펋l��&t�f���t�����     8D�     �aig���^\�ZI�bRl��b}9�    p��    �C�t���^^�Zm�v�E�a��{� t    �!3p    �wk��2;}y�$i�b��-���oCw     :w     ~�$I�l��t��-�r��ߟ�ZM�    ���    �$�'�//Ӵ��1)����Ҹ    �S1p    �W%I�>���L�a�bRU�����E�T�[     >�     ���9�<��vF��%���ur�v    �O�:     �x���y��eE��I]��r�ꢩ�i�    �c�U     ~�(��}�7[��M���ϛ��    �g`�    �����Bw@\�$_�>����    �X�    �O���ht��qi����yU���K     ���;     ��?x��Ə�; 6���}���     8v�     �Z�V�۟��ٓ�; 6w����r�    �>0p    ���e�l��&t�f���tW�OBw     ��     �\�;.��s�v�����l[����     �O�    3�Nf/�Z��	�1Y�/'��z�    �1p    ���i�̌��_��I���i�    ����    �J���d��e;I��-��n>Z�?=�    p_�    �3I�V��7��v�
�1)w�`���Q�    ����    �I���f/�Ҵ��1)˻~�x{�j5I�    ����    ��H��鳫Ng�]1��׽����V�6n    ��    �^H����n�d�bRU�N>}�4�;    �8�    ���'7��d�bR7�4���h�*�    �3p    8r��/����u��I�����u]vB�     ���    �����`��.tĤi�v~��y]�[     �g�     Gj0:[�F���&Y.^�WU�]    ��2p    8B���|4�j���$���YU���K     �e�     G�۟��ٓ�; 6���̇�;     ���    �H��m�����; 6w����r�    �_g�    p$��h�͞]�ZI�b���v�+�'�;     �m�     G M�l���j��?X��Ͷ��I�     ~w    ��N{ev�򪝤u��I��Ί��4t     ���;    �k�;U6}y�N:U��IQ|���=�    �c�    p��$���7�i�ۇn��lw��u���     �q�     (I�����e����-�r�V�v    �Ce�    pp��d����B�@L��U?_�=o��$t     ��    �$����u���K &�����ߜ�Z�q;    �3p    8 ������t�bRU�N>}�4�{    ��    �@Əo������;��8�>\�==��7����"���%&N�c43=KOW=/��q�Ւ��X#��9fΑ�IJ]�~�������     ~?�;    �%0��|>����������OR�F��     �v�    n2��z��������j��ORlJo    ���    �xzs�X�����/^<������K     x��     ՌW�r��ץw���~����k'��     ��	�    �n�Ս{�.��f}��n=+�    �wC�    00�hv�q��Y1��C�Y?��;\�K�     ���    H]O�+q;��v���q���     �-�;    �@TUsZ�:V�:��C�n��y�����     �=�;    � Tը_ݼ��*���[`H��W�}�Ս�;     x?�     ��X�������������E����w     ���    ��yy��t������������    ��%p    (&��Ͼj����n_<�    \Cw    �B7�����]�0$�i;Y�x�q9��    ��'p    (`���ד�Ͷ��өo���    �3�;    �{6[��v:�`SzI�G��>ι��    �sH    �M����?�(��$���x�������     ��    �'��������C�r_]<�INݨ�     ��    ����v���M�0$9�j��ORhJo    `�     �XӬv����.��%ǋ�>�����     �C�    ���b��y��;`Xr\?�Q�m���     0,w    �w����Ս{_�s�-0$����6��;     �;    �;P��nu��Y�Tz�v���x1/�    �a�    �e1������*���[`H�맷�o��w     0\w    ��(�:���˿�z|*�������a���;     6�;    �[c�V7?�W]O��[`H��W�}����w     0|w    ��"�卻�F��������E����w     p9�J     �
g�^ԣeL9Lb9Ęb9�b)�Ko���p|1k����     .�;    ��4[��ԣ9�0������r�1�B�!��r~��ë��1�E�\Z�q=ݾ���;     �\�     ��t����~�'�C�!�P�����1� �!�����A|!���c1��C��ˋ����鴝l.��(���    �5�;    �o4�}�O>:���B!��� ���W�����琫*��s�1�c�!�r9�w�B��C�~������     ��;    �o�L?�Of���w|�?n���~|3|!��
BL߅�!�\Ő��o����ŷ�D�    �o%p    ������w�w�6?u+|���Wm|!�C�!��VH!�s�1f<?��^?�I�}]z     ���    �W57�����?��
�/��9T�#�7�b��&�������&��B9��B�_)��ŷ�$��s     ~�     �P�,���������˜�!����e��'�*Ɣcz���ݯ)��b����m�9U�o|��cSz     ���    ����i�<߈��RU�U��e�C9�S�!��>�C1�B
�K ǋ�>�����     ��;    �Ϩ�I??;߄X��r��r�r����|9���)��b�)���f^�q���G}���^    ��!p    ��j��gY�8S�o9�B�� ��1�r!�R����R��s�_|�u�Y�     \-w    ���&��؈�'��Crr��_�9Ƙ���n~!�B���^=�����_,J�     ���    �7�΋����&��~�cΡ�C�x�{!�cHU)�c�B
9����/o�߬J�     �j�    �H�g�몞	���BUΡzy�{���c�1�sH!�cH1�cN9�����?o�w_�(�    ��K�    �1�W�6u��K/�=�!��Br|�B�9�ؿ��S�1�1\��}��j�o�u��     �6�;    �f��6���Tz�c�9�^��ի^��}��f�n��C�     \}w    �W��;�f|�+��K�����Y����    �� p    !L�lǓ��wpE���=�cz��C�C�)�a���q=ݼ��r,�    ��A�    \{����d�ɡ���BUΡ�oF����bc�c�r
9�bSCݩo.��     �_w    �Zk&&�O��wp��s����e�C�!�R��y���������G��W?��     ���   �kk4�y�-w��C�9�9�:�q�{�bCJ!�������{J]}����s���5    ���    �Rݬ����6�Xz
�
1����������c�c�U����_��S>��|��I�    @w    �کG�n�:߈۹2r�9���k�_��C�1���[�c�c�駾D�}����ǩ?6�e3     �w    �Z���i����v��bΡ�!���y����͛�s\�x�q���E7    p�	�   �k��'����&�W]�u���]?Z�]+n    ����?    ��U��sq;�@����ԭ��     ��    ��b���몚��S`8r�m��O�q;     �!p    ��*/�z*n�7�Og��I�     �&�;    p�Uy��|S����}�t�����     �I�    \Q1�Ww7�fu*���69�    $�;    p%͖�mF�q;��x����>���     ?E�    \9�ş�f|�+����7����w     ��"p    ������d�ѡ��Sw1ڭ/K�     ��#p    ��f��~2��/����u+n    ���    WB3��0��iWzI��z���*�Ko    �_B�    \z���q��Ӗ�C��}�]?\�Ћ�    �4�    ��V7�n���A��I�P�뇫�N�     p�8�    .������^K���ŃeJG�      �tn    �RUO����&Dǜ�O��x�J�X��     ��'?    ��SU�4?���q�Ko��H��x�L�^�    ��%p    .��j�����������v�h����     �=�    ���<_���j�JO��ȡ]?^�ݺ)�     ~/�;    pITyqv��ꙸ���n�d~�^�K/    ��A�    \U��>����/��d�}:��LJ�     ��E�    �l��vԬN�w���/���i�     �6	�   �A�.�l��fWz�a�lr��kVz     �mw    `�&�?��ɇ��;`H���Ǉ���     x�    � Mf�w��Ǉ�;`H��y��>Y��     ��    �f��a2�t_zɩ��֏��w     ��$p    e4�y�-w����M݊�    ��    �`�ͪ�/�nC����`�}[o/�BH�     \yw    `�f�-V�q;���}ծ.C�1     ��    @qU=;���R>�v�p���Y>     ׆Cq    ��������Jx-�.�/��J��    ���`    (���i~�/�*6����O��x�J�X��     ��    (#�y�:����^<\�~/n    �Z�    �yqv���i*��#���Ѳ��Q�%     P��    xϪ<?����E_z	G�����M�%     P��    x�b���mF�թ��v�'���Ÿ�     (M�    �7��g�Qs&n�7�ڧ���ͤ�     �;    �^Ln����C��i��jZz     ��    x�&�Ow��G��;`H�g������;     `H�    �;5�~���n�K�!9�ڧ��;     `h�    �;�L>8L���N��f�}�(�     �H�    �����lq�-����]����v     �	w    ୫�U7_�݆KO����mݮ/CH�     ��    �[U���b��F������W�v     ���    �[S��~vv�	��#|'��j�~���    ���	    x+�j��g��U��[`(R>�v�`�S�<     ~�    ��VUͫ����+)w��x�J�v     ���    �O��|u]U�Tz
E��q{�Ko    ��D�    �U^����z*n���оx�L�^�     ���    ���<_}���E_z	G���e߷��K     �2�    ��|��vԬN�w�p��n���uSz	     \Vw    �W�-�nF�ͮ��vۿ�O����K     �2�    ��d������v��Yw�zRz     \vw    ���>�M�J�!9��1��_MK�     ��@�    �"���dv{_z�a�lr��sVz     \w    �g5�[���O��;`H���Ǉ���    �n�    IDAT �J�    ��4jng���b�)0]���o�,J�     ��F�    ��z���{[q;�v�֣��q;     �w    ࿪��iqv���k}�����e�     ��;    �#U=��g�o!�k�o�틇+q;     �;�N    ?PU�4?�˺�M.��"��j�~���    �;$p    �WUM�����R>�v�p�S�L     �1��    �+u����U5I���P����ŃUJG��     �8�    BU^�}��ꙸ^��ۋ��u�-     p]�   �ڋa����G˾��ڋǋ����     �	�   ����>ی��S�09l���iӔ^     ׍�    ����ζinu�w�p�Ю��軵�     
�   �55�}�O><��Ñ�n����{>.�     �+�;    \C����dv{_zɮ�r�����     י�    ��f��a2�T�o8��1��Ϧ�w     �u'p   �kd4�y�-w����&��?g�w      w    �6�f�͗w�!��S`0��oƇ���     �%�;    \�h�-V�q;�v�.F��E�     �kw    ��z��W���o�O��]?^��KO     � p   �+���i~v�H������^<Z����     �;    \Q�j��������^I���^<\�Ћ�    `��    p�:/V��U5I���P�t����U��v     *�;    \9U^��_W�T��������2�ι8     ��|    �R�<_}���y_z	Eʧ�^<X�t�Ko     �7�;    \!���ͨY�J��H��x�L�^�     ���    �����f�����rخ-SߎJ/     ~�;    \�ş�f|�+��#�v�x�w��     ���   �%7�}�O>:��Ñ�n�d~�^�K/     ~�;    \b����dv{_zɮ}:��LJ�      ~=�;    \R��������;`Hv��Y��jZz     ���   �57�����!��S`0�g�n�L�     ���    .��Yv�ս��^;�ڧ��;     ��G�    �H]�O���F��u��f�}�(�     ���    pIT�����oBt��9u�����     ���$    .�����_�1�r�-0}��[q;     \)w    �X5i~v]�F������/�BH��     ���   ���:/V�몚��S`(R�����zq;     \1w    �*/���U=��+)�v�p����6     \A     � Uy��|S׋������^<X�tt�     W��     0@���mG��TzEΧ�^<X�t�Ko     ��;    �tqgیou�w�p��^<\�~/n    �+N�    2���O><��Ñ�v�h����     ���   �@Lf�w��'��;`8rh׏}�nJ/     ��;    @3��0�}�/��#�����Խ�^     �?w    (��<�w��;`Hvۧ���ͤ�     ���   @Au��f˻�b�)0���iw�jZz     ��	�   ���Yv���F����&���f�w      e�   �������{nn�7_���y�     @9w    xϪz�/��ob��[`(��y��>Y��     �%p   �����4_������b�[?^��     �'p   ��%�y�����I*=��?m�V�     �"p   ����˳�몞��ᕾo��ţU)��     ��    ޹*�W�o�zޗ^C��}ծ.C���     ���    �N�0_�݌�թ�����]?X�trF     ���    �͖�mF�q;��r�]��9�     ~�    xG&�?���VWzEΧ�^<X�t�Ko     �I�    ��d��n2��PzG
���e���v     �'	�   �-O?�Of���w�p�]?Z�};*�     6�;    �E���t��]�09��ǋ�[7��      �'p   ��d��<�w��;`8r�m��O���K     ��A�    oA�,����6�Xz
Ʈ}:��LJ�      .�;    �NU=?-��q;�v��c����     \.w    ��z�/��7!:j����&��?g�w      ���n    �U�8���c��[`(���Ǉ���     �r�   �oPUM���_W���+��y��>Y��     \^w    ��b���uUMR�)0��bԮ��     ���    ~�*/���U=��+}�����e)��     \nw    �Ū<_}���E_z	E��z{�p%n     ��;    �B��g�Q�:��C��}�]?Z�܋�    ��B�    ��tqg;jnv�w�P�|����*��93     ��x�     ?c2�S;�|x,��"�.�/���     x�<|    ��a2���L?>��C��)�V)��[     ��G�    ?��|p��>ݗ�ÑC���2�{q;     �N�   ��og�;m�09l��}ߎJ/     �.�;    ��Qs�8_�݆KO��ȡ��m�w��     �j�   ��f��W����vۿ�O����K     ��O�    �T���X�o���ڮ�r�����     \w    !Tդ��}�qd�v��v�g��;     ����:    ������������[`(�g���;     ��E�   ��VUM��������Ǉ���     ���   p��y�����I*����7��E�     ��$p   ������ަ�}�%0�n=ڭ��     ��   ��b���mF�թ��������2�Ko     �/�;    ��l��fԜ���Է���Õ�     (M�   ��2]��6�[]�0��W/on���     @qw    ������x�������]?\��9+     �C    �����n2��/��"�.�/�R::'     Ã    ��f��a2�T���p��ŃUJ���     �7	�   �Қ���lq�-��#����"�{q;     08w    ���Yu���m��������iJ/     �o�    \Iu=?-V�o������}��     �%p   �ʩ�i?;;�8������}~ꞏK/     �_<�   �J��q���_Wq�Ko��ص_κ�ד�;      ~��   �+���Wq{#n�W�N���i�      ���   ��!�y�����I*=��x�����Ǭ�     �_J�   �P��������vx�;~��_��     �k�   ��<_}���E_z	ũ��6_,K�      ���    \j����Y�J�O��]?^��KO     ���    \Z���ͨ�ѕ�C���z{�hB���      �w    .����m3�%n�WR�����e��     ���    \:�٧����C�0)�v�`��ə/     p�y�   ���L?�Of���w�P������2��y/     p�y�   ���Lnf�?�JH�ۋ���u�-      o��   �Ka��8���!��S` Rh/.S��     W��   ����e7_�ۊ��;9l׏��oG��      �Mw    �����|#n���Ю/�nݔ^     �	�   �������7���;9�O��Ÿ�     �w��A    ���i~��u�\zŮ}:��LJ�      xW�    N��4?�/n�7�ۧ�n�մ�     �wI�   ���y�:_W�$�^Cq�?�����     ��'p   `@��8�|]�3q;�r<|=>�O�w      �w �c�  �B�սM=Z����Pt��f�}�(� �m���|   �Y ��+��RhR�u�)  �0[}�5g��;`(N��h�~�,� �mI)6}��1�t   �iw ສ�>�S�� �Lw�Ms�+����u+n ���¨��2�Д�   �� �^b9�ѩM��-A  0���O><��C���޾x�
!�� ��r�}_�R���   ?4*=  �=��>���  �1���M��JH��ڮ.C��� \y)UM�yT�as>��   ���k���  ��L>8Lf��KH�P�뇫�N�m��#�؟�<�j��   7� W^�}��v ���og�;m�0)w��x�L�(n ���>��Gu��1��  �5�a	 p5�r
�S���v �a��U7_��ߦA!��O��x�J�X�� PT�U��y
�4��   �-�; p��Ǧ�A 00�h�-V�q;|'����2�{?�  �B�!�aܧjB�=   \Cw �J�9�}�M���9  S��~����v�^���e߷��K  �&�P����9L=�  ��Ń ઈ)��˰=�� ���q���_�8���Bȡ]?^�ݺ)� `�b�Sǐꪊ��s*�   x��]w ��sk; ��ŪI���*6�v!���n�d~�^�K/ �r�꾏��ä�   ��s�; pi�b��(���v ���u^�j�Exe�>�u�o�Y  �F1�j��4����9�   �(�� �UuJ�y� 0LU^��_W�Tx�v��v������{��4����[���>UU�cQ�P�H$g�@H`%��|���Er�H� �� ��شE� 5$�D�C�4�"(���(6�p`�!�(pDٖ(rf�{�gzM���յ�Z��gHΡU���y����z��}�{��;  �խ�ܻ��o�   ��0 `���y��֚Z�  �F�:�z�^7���%�(�����_���  Xz5R�iZjL#%��  `�[  ܹ�r�}�� ���m�{o�o�[w���y������u �*)��K�����Տk  `E8� X
��`��ȸ `�M7߽7��f����\���l��  XI5��c��4n�   �w `ѥR��śg  ��d�G��'�;`Q�Ov����7[w  ����q��F$��  `ٹ� Y�K���� ���w��?xܺE���� �M-1��n�F�[�    ��X X8]��5��}��Z�  ��F�:O<j��"���Υ��� �<�H9�i�1M��e   XF��  ��"��\� �H?�cǓ���EQ�Qw�{q3"�� h���/���8�Zs�   ��9� X��`^�� �L���nN7~� |����(�f:�}j���{�  �����Qj�N   , @s]JQJ��İ�j �$���l�=���pK�'�`穭RN�w X)JI�R�YJ��   ,Z �ֺ��R}/ X&��l����q;�R��ָ=Z�  ��J��IN�5Rߺ   xs�d @)���s�Nm X.�`�gދ���R�`��f�G��  ��F�9MK�iJ~�   �j�:  XK)��k�  `�tݨ�.<��Ұ�n��Pc��f�� ,�R��Ft]*G)"��   ��c� �sUkrI��  K(u}�]xd�K�q;DDD�����d�o] �ݩ%�t�1j�   |7w �|��Zb�Kk���  �&���û]7.�S`1�8�v6?�a ��j���I�1Mɡ,   �(���JN}�1h ����ƅ�w��Ըn;<�:=9~yܺ ��WJן��6   ,w ���.�ԗZ}�  XJ]�m�wo0�ȭK`Q�099�֤u  ���n^�Y�ԷN  �ugh ��Qk���V�v XRӭ��[���(�����_���  ��H9�i�1���  ��a�  `%���Щ�  �m���~߿��u,���/����Zw  p�J���Eץr�"��
   Ι� p�R�K�� ��x����;n��E1?���_�h� ���%��Y�Էn  �ucx ��Qk���V�n Xb�郇��?n��b~�3<�}Ƹ `�ԔrN�Rc)��  �sb� ܷ�JN}.1h� ����?p<���u,�����7#�A ��*��s�f�<_  ��� �_ݼ����{ ���Go�9�x�u,���;��� �%��m�H}�   Xu�h ��I��p����{  ,�A�u2�|�~��vQ�Q��{i3j�G �-5R�iZ����'   83� �]K������-  ܿA�y����}�R��t�{q���O �>9�(ט��y;   �� ����%�R��  +�L���8�n+�$�xj����y  xC�t�����Ұu   �i �;Vk�9�Z��  VA7���4��[`Ԙ�����J9��*  �R���<f�Ƥu   �w �-u)���s	'�  ����مGv���U5n\�,�ȸ ���"�n�K�"%��   �)0p �J:�1*�7  ��4����w�42n������{q3�}?� �����9m�?�  ��d� ��.���N� X]ݸ��n7���%�j�=��Ov��%  ,�].iV#|�  ��`� ��Z�`����� ���ζ޻7l��%�j�?;�߼>j] ���)圦�Ƥu
   ,+w ໥�R�ϥ[�  p�R̶޳7��K`Q<?=9~yܺ �U�"�n�k�"%��   �]2p ��)��R}G  X5���������&'Gל�	 �����sڈ�A�   X&�k �m����k��  ���Ə��NZw��8>�6>>|qں �5P���nV#F�S   `Y� QK���V�v �3���p4�����(n�<:>�:k� ���r�&5��'�   ��\>��R�R����Q VQ?���������(NN��G�W6Zw  ��r�QɱɛT  �����J��I��R}  XE�����w��E1?��>c� @S�t�y�6"��g   ����5�}�N� XE���oN7:h��"�����͈� ��jt�f5b�:   ��; ��Zc�Kk��  +h�o��6߽~�Q��`���-�v  J��s7��MZ�   ��1p�u�R�}.ᵧ  +�������-%u�Nn��(  XH9�(�n)��
   ���H)�:*�g? �����q��H��ADD�7���ŭRN�Q  ��j��<�FM.�    �� �A7/���O �U�u�2���nJ�ںA��t���V)7�� `9�ԕ�6jİu
   �� ��Zc0���  ����2���n�z�v�[����'�J>�n ��Qk��ӬF�n  ���`E��\�� ��Ҡζ��qi������卒��� XR)rN�ݤu	   �b� �&�(%�\  `�uu��û�`j�Qc��f����K  �~��\�Y���   �w X!)"�\G��� Xm]�m�wo0�ȭK`1�8ܿ2�'���  ��Zb8ϱQSr�  ���B VG7/��Ns Xq����[���(��NO��3n�  �����Q#��S   ���
�5�l� ������o?i���������[��  pVj��s��H��-   p�`���\�� �Ƴw������k㓣k��  ��9�I�n�)?   �Υ/ ,�����s�A�  ��x���x�Cǭ;`Q�<������u  ���c�s7����  ��e� K(E���T��  ����x�Σ��(NN��G��n��  �j��<�FM�3   V�^ X>ݼD_k8� `Go�9�x�a�X�������  �TM]αQ#y�+   +�� �K�K� ��a�����wy�780n �[jJ��Y�ԷN  ��d� K���s��V�& �50n�̶�c���?�߹�Q�Q  ��j��cZj�N  ��b��dC�    IDAT K�����  ��n0�o\xxϸn)��;ؽ���Q  ��IQJ���%   p�`�u)���s�A�  �G׍���{�ܶ�[J9�v�ڪe�  �D�]�k7��  `�y( �*������  k��Fe����R_[��"(�$�<�Yʉ�"  ���0�n���ü���/_h�  �ƃ! XL)�:*��� X]חمG���R��`穭Rnz�  ܅Zb0�i�����ã��'�3�Ժ  V�Z X8)�}�NW X�:�z�^׍K�X%v.n�|d�  �����)�Ng쥗��/����;  `���b�� �MWg޳�f�u	,����6K>�. �eVk�yN��o���&�|���_i�  ��� D�1���k���  k#�l�={��ּu	,���7�ɮ  ��)瘖�ƭS`��x����?���u	  �w X ��0�p:! ���n��ް�`�Q�p��l~rcԺ  VK�RҸD7i]���O\����}���Z�  ��3p���Qr��Ġu  �k���~?z�u,�Ã�ӓ��8U  �H�1ʵ�E�7������Փ��|�o��t�  Xf� �JJ1ϩ/>� ��x�����7[w��8:�:=9���$ ����\�Y$#w8+7O�������|���Z�  ��2��6R�uTj�Y �f�����Zw��8>�6�yt͸  �I-1��n#�� ������k�'_�޾�`�  XF.X���H)��ku:
 ����?p<��Ӹn�y������u  ���<���4h��jg0�Ʒ6���]��[  `��������  k����t㡃��(Nn���_�h�  k��4/i���ʷ���.��]l�  ��� �O�K�Z�� �̠�:�n�{?��""b~�3<�{z�u  ��i�Ӭ��i8#Ͻ0y�/b��m�  ��� �A�1���� ��`�y����q;ܒ���`��q;  ,�)�cV#F�S`U]�2�w��s�7Zw  ���+l 8c�� ���:R�nPO�_�Q��S�� XL���l����RO�����n0*�[ �jN��8�R��c�u5u)�[������ɋ�������ŗ?���[�  ��3��3TKs�A��������;N��ƅw�l���O�� X]���֏��  �8>|qr|�´u�FR��Ʃ+)�8j]�&׈�?1��'������?n�  ��		 pF��    �e�K7*����Ut�K_���ß��K�n �Ef� �-EԚ��    ��TJ�r�Y�H�[`���O<����f�n �Ee� ��K%G�K5n     �V�ݰ�n����Խ|�����{O��  �Ee� �%E�s�K��
     ,�Rb8/1K)��){��䡿����i�  ��  NG�9F�V��     �ʨ����0r���ԕ��>���߷�  �Ec� �/�}�^�	     ������6jJ6p�jJ��Kӿ�������-  �H\|�}H���    ��W��96"Ҡu
����_]��g>�}�[  `Q�������     ���)�K�E2r��tt��vy���_��h�  ��� �M�K�Z��    ��Q#�s����)�Jv��'�p;  `���3n     �W��s7�)��)z������?l�  ����1n     ��rN�F�p���:��m����  В�; ܱ��s���      q{��ѷN���R|����|��|�u
  �b� w$u�\ݜ     �.)n����%�*�%�'���_���O�n ���-�����      o$E�ib����8������K_zq�u  �7w x5�h����      o�Ց{�\N�+��������  p������$"�N     X)r�I�1n]��������~�u  �'w x��8���W     �����nl���ɧ�������[w  �y1p��Qj�v     �{VJ7�5&�;`Ԛ������;�u  �w x�1)%�     ܧ\���;����.}���lo_{�u  �5w ��D7)���      X�t�F�p����oo|�u  �5w �W��a�     p�J�F�vF�p
^ze������o�  g����WjL��     �N)a����s�?����u  �w �Z�ݤ��o�     ��n�����S��'.M��c����o�  g����uk���v     ��RJg���$G��˛�㧾��C�[  ����j�v     �J�F%���~���.��e�  8m� ��Rc�Kg�     �H�ݨ�4n����+������N�  8M� ��1)��      ͕�ƥ��;ܧ���ԣ���\�  8-� ��RӸd�v     �EQJg���F�^?�����S�[  �4��J�q)^s	     �h�����tݥ�7~k{���[  �~���n��;7E     T)i\#y/܇��������  ��e��J��F��      �.E�11r����K���O����  p?�XY5b�sLZw      p'^���;ܳO\��G�~v�íK  �^���n���$"�N     ����9Mj��u	,�\#�~���?����u  �w V�q;     �2K�sL����w�o<3�����u  �-w VJ���     ���;ܯ���W�~�u  �-w V��q�Ը     `����j�G���[}���j�  w����P#��tNn     X))rN�a����O<=���~���[�  ��2p`��H�\�iT�v     ��S#��M#Ҡu
,�㓮����omoW? `)���j� ���     ��i^bVS�s�{���p���޿h�  w K+�t봎���     V]M)�4�����3�O~���7~�u  �} ,��R:�i#��2     ��Q��9�"y�/ܭO>=�k�����n �7c��I)�K��     ����\�Y$o���u|�uO]���?��uܺ  ވa  �%Eʥ�j�A�      ڨ%�T'��=��3���{�ߺ  ވ�; ˣ�ȥ����     ��Z�A�1m����s���ۻ�m�  x=� ,�2例İu      ���nX��;ܭO^��G�֟j�  �����P���}�      K)]_j7i���xޥK�l�֗���F�  x-w ^�1)9F�;      XL�Ĩ���es}o8��6~�u  ���; �F���     �J��F�p���:�����/��  �W���j�(��:I      �H)i\Û��nԈx���C������n �w TMi�s�D��)      ,�9�IMiغ���I����ֺ  "�X@5� �45n     ���9M#�A�X&߾1���'w�Һ  �X,)�\bպ     �{T#�s�"�E�ݸ�����=~��;  Xo.� X)�4�i5�     pjJ���R��	�T.)���䗷���u  ����Ő"�K�EM>�      85�yI�o�;�4^����Zw  ���X�t�Z�A�      VK-1ȵ���er���]?���?��  `=��\�ݤ���      `5��RcҺ�G��.���G����. `���T�1.%F�;      Xm�t�Rcܺ��I�ҥK��u{�:� �se�@35R_Jr     �sQJ׈�u,�����ý޺ ��b�@5b�K�D��)      ���t�iк����&�c�����  �w �]�䒦Q��     8g5R.1�)�L���G�۟����n `=�X�|��r�Q�q;      mԔr�Y$2��88�W�L���  �w �MJ�rI��>      h��.�n����<��������׺ ��g`���"楛���)      QK楛���P�˓?��_��S�K  Xm� ���cZK[w      �k��R�����KO<3���  �6w �\�1.��[w      ��)��K�q�X�~e��|j�� �3c����})��@      Z)i\#y#1܁KW�����?i� �j2p��A.�$"�     ���"��FĠu	,�yI���㿷�]�( �Sg���H)�K�F�n     `IԔ楛F�����~������  `��p�R�\�,��      �L�.�nf�o����=���|�u  ����SWJLj��F      �S-1(%&�;`������_���_�u  ����SUj�K���      p?J��Rcܺ���p����u  ����SSS����     `%���5�a�XtW�?���Ϸ�  `5�pJ� �4�H�C      ����9�1h]��FēW��޾�`�  ���; �/E��4�j�     ���)�K7M)yob��^ޙ�n�  ���; �'E�%fQ}�      ��jt�f�u�𦮾4~����|�u  ����RJLj鼒     ��VKJ�I�Xd5"����c�o��p�  ���; �������;      �<����Ƹu,���n�ͯׯ��  `y�pOjJ�R��w      ��RҸ�4l���ʋ�w��/���  ,'w �Z�䜦�u
      ��9�i��.�EU#�+ӏo�Z}G�  ���; w'Eʥ�F�n     `M����R������`��S��ۺ ��c��]�%�Q}~      ��jt9�i�Xd�>?}�G>{c�u  ��@�;V"&�t��      �j톥Ƹu,���|��~���-  ,w �HMiXr��      �ERJהo`�>�����  `y���Rt9�iDj]      &E�1�d�o��F�<���?ֺ ����
�7�R�\�iT�v      x]5�z���(x]%R����/~�ׯ?к ��g����%&�Ġu      ,�ZbPjLZw���?/��૭;  X|� ��Rc\J׷�      �ePJ��H�����~q��~���u  �����U#J��|     ���sL"%oH�בK��g'�Һ ��f���K)Ւ�Q#�N     ��b�c)y�����p�W?��ۭ;  X\� |�."�:+�g      ܓ�R.i����W�������m� �br)�w)����ye"      ܇ZbPJLZw�"�9O�ꋣԺ ��d���V#�%Ǩu      ����Q�Է�E��˓>򙝿ݺ ��c�@DDԈA.�	      p�n?��e�>5�yy�_|��/?Ժ ��b�@DJ)�n5R�      X)5Ҽ�i��Y|���������ٺ ��b�@�\�Q}&      ����+ަ�빗f?���]�T�  �1#��+5Ƶv��      ��J��F��ES#���O�K/n�n `1���4(�s      �A.i��;`���'�����  ,w�5�R�yIӨ�Z�      �Z���%�)yF��F��'��ӭ;  h��`M���>      �\����MZg����.^���  �g���j�Q)]ߺ      �Q��׈Q�X4/_m}��7�~�  �2pX?�\Ҹu      ��\�qM�n����&?��_�{�u  �PX#)E��4��u      ����4������q7������  �c��Fr�IT�@      �"�%�t޾��ʋ�G�ܷ�|�  �0rX5R_J׷�       ��ĨF�^��..=7���  �a��Rt�Ĥu      ��r�IM������~�C�7~�u  �����K�r�QSj�      ���R)i���k<���?����m� ��2pXq�t�Zbк      xc�ĠD�[w�"9>t�<7�g�;  8_� +�F��Ĩu      ��JN�iغɳ�O���^�˭;  8?� �*E�K7i�      ܩ�Ĵ&{xU��g�N~�u  ����ʥ�F�Ժ      �5�Zb�:�����C�;��u  ���`��ƵĠu      p�J��Ƹu,�����?�ŗn� ��3pX9iP��]      ��J�FɡVp��I�=m럶�  �����4/i�Zw       ��F�5M"y��z���?��o��;  8[� +��n���      �
j�A����*5��g��ں ��e	�"jJ�R�u      pzJN�1l������[����Zw  pv�V@J)���vB      X1)j�&�<�W=�\��~����  �w��K�DMnh     �
*5�RbҺ���`�����v�  Ά�;����R��u      pvJ���sA�����?��^���  �>w�%VSt�t��      ���%Mj������ܥ^���  �>= K���F�Ժ      85R)ݤu,�������\��[w  p���T�1����       �O-1,5��"�D�+/��ܺ ��e���jĠ�nԺ      8��:"�;;�Ƈ�o���  �w�e�"��M�Fj�      4P#��M"<3����W�v{���;  8� K����4      Xg�ĠD�[w�"88�?��v�  N��;��)���Q�      ���ӨFr8Dĳ���{���d�  ;��H9wo      nI�K�F�n�Sz�Z��[w  p���D�n���      �k��j�q�XW�������3�;  �?�� � �A�u�:      X<��QD���JM��3��Zw  p�]��K���
      �+E�i*B\{y�����o� ��3pXp�ĸ�p�      ��j�A��АR\~��x�  ;�BK�R��P      �[*�E8<���ӿ�}�j� ��1pX`�^#�-�      ���r�&�3`\~n��>��uܺ ��g���J�q-NW       �\-1(5�zY{{�ݰ|u�k� ��3pX@5����      �J��(�M\~�����+{��  �X@��i�H�;      �%T#��M[g@k�']��g�[w  pw�L�1�%�;      ��UKj$o�f�=���'��|�'[w������Y�����Z紵)�h)�)
HH�RH��XP4�@Jh�=�ª��S
��^h�)&�7���1å�s����e���/'��e��c������/��1��  <8w�]�1�2      �jy�´�o������9  xp>b vȪ�Q��s       #P��6���}���-��'�� ����#*rY-�s       �Q-��i&�*���a�v�  <w�Pê�A�      ����p��^�fҞ����}��O�� ��Sp�m5F9P      6�"W�{ǀ�*2�����s  ���:��yU�{�       ƫ�aQ��%��+W����/_�w  ^��;@_�jiR      �q�UF���������� �W���QUDY�     �-�Z�e��ӕ��|�����9  xyJ� �T�l��      آV��L}&�O�^��w  ^��NZ�ax�      ئ�l-{ǀ����y�/��v�  �4w�*bYm���      LO��W�w�鏾����  xi
� ۖ����c       ӵjq���f�Nnϖ?ut�ӽs  �g)�lYUD9(      :��Vs1m�<:�y�  |)w����jU��)       ڪ�9�z�y:[\���� �/���E�����     �]���:�z���~���[y�  `�(�lI�8��       ;��0��P3Y���|��O�K�  �
� ې���B      ��Y�<��5�����m�;y�(    IDAT ��Pp؂���(B      �����w����a^���3�s  �w���y�X��      �rZ�EE�{�^>������ ����I�Z�t       캌VÁ&	Su��l~�����s  ���Q��2*��      �Ϋ�����9���}�{tT�� :�!ؔ�l5,{�       xP��eff����;������� `��6��p~      ��Q��JSܙ��>u��3  L��;�F�l�j�;      ��j�ZFĬw����|�S�p��z�  �2w�XU���      �^�h5���d}���� `��֬"��      ���Z�+s�;�pr{��飓�; �T)��W��I      ��[��0���L�瞞�X�  S���F�bem      F�bh-��c@�O�?}t�7z�  �"%L�u��V��      `4Z��4ŝI�³��w �)RpX���0��|      ��T��w���٣?�� `j��"g��w
      �uk�ZFĬw��s��� `j�֠U���      �(e�Lqg��\[��C��#�s  L��;�U䢵��      `�Z�ye�{�m��x���'{�  �w����UK�
      ��[��0���L�ӗ_������; �T(�\@k����      P1���1`�V-���ӽs  L�R&�yef���      0��ef����<���_��'�z{�  S��pN��A���      �	��U�A��mg���7^��{�  �w���ZŢw      �mkmXT�0=�}z��GGW�\�  c�c��j0�      ����6�����=��ޝ�~�  c���*b֪Lo      &k�jQ��9`۾p��;��j�; ��)�<�V�A�      LZFհ����a~�n�n�  c���02g��/�     ��k-�i�;��gf?�; ��)�<�U���       vEk��ɹ~2?��/]�H�  c����*r^-L       �S����
6��ԥ����  0V
� �U��       �kZs���\�r��>q�z�  #w�PK��      ��j1��E��M׮�o�� 0F
� �.WmX�      ��V-�P��/^���?]o� `l|Z ��V���^      ��ʡZƤ��������; ��(l����V�      �U�s/cg��M_|z�7zg  w�W�j��J0       ��U�LqgZn���?}t�7z�  w������      <�V�2�w���K?�; ��(���U��(/       �"[���1`�._^��O]��s  ���;�K��Vâw      �}�jXd�abLFEƟ|q��9  �B��%�2�      �\*rUe�;���僯��_��s  ���;��df�fz;      �y�6,�w&�~�|���?�� 0
� /Қ��       R��Ųwئ/>�������� ���^(#W���      \P�\��Δܹ;̮���w �}����� �      ��Udke�;�������  ���������      �Iհ�CƘ����{�ɫ��; �>Sp�S��2��
      ��TE�Z���dTT<ue�k�s  �3w��禷�C      �uk���3)O_Z��S�z�5�s  �+w�x~z{:P      X�JSܙ��g�����]�  �J� "��a
      �����dc2��r�=�3  �+w`�ZŲ�A
      ��Tf+Sܙ�k'�G?��g�Q�  �H�����fz;      �Ƶ�e��cLDf|��#O� ��܁I[�XF�      �M�̪\���쥃�::z�M�s  �w`�Lo      آU3ŝ�8[���#�� `�(�����v      ���LqgJ������3  �w`���V�C      �-[���6�q|k~��'���w �}��LR�XFY      ��r�ɘ�K��?�; �>Q�&��v      �~Z���t<{e�棣g��w �}��LNeΫŬw      ���6�"ӽ-�p�����w �}��LNki       @g���3��<}y��3  �w`jf�j�;      ��U�ye�0	ׯ���'���; �>� LJ�XFd�       DFy�����x���+�s  �w`223[��      �V��4��ix���GG^� x5
��d�VQF       vFE6Sܙ�ӻ��Z�Z�  �N�����U��9       �RU�LSܙ�KW�� `�)���j�4�      `�TE�J˘��������{�  �e
��$4��      v֪�w؆U˸r��w{�  �e
���U�"�z      ��*�ʜ���������  ��>��k��       ���<���ƭ����8���9  v��;0j1���9       xe�b��w�����c�3  �*w`�Z���       {�5/t3�^9|��� `)��U�C����      ��i���,��ݳ��]���9  v�`��r��c       ��2�y��i�r���{g  �E
��Xek��      ����\D�f��]��x������9  v��;0J��J       ��2�r�;l��*����z�  �5
��(�Lo      �S�j�;l�3�f��; ��QpF�"g�b�;       �Sm�E�{_F����}��7�� �K܁�)��      �{���e��"._����9  v��;0*����y�       \L�a�;lڳ��w �]���ʪ�2�      �ޫ���wF�����#�|���9  v��;0*��E�       ��;`&!3���O� �+܁Ѩ�y�u      `4*�ʜ���v���/��  �+A��h���      ��*w��ޭ���瞼���9  v��;0C��}      ����y���������  v��?0
�b��c       �vUa�;�w���m�3  �w`�ed�a�;       ��Z."M=c�N�͆���� �7w`�UŢ�A      �hUfU�{ǀM�|<���  zSp�^�0�      `�j�;lڥ����  Л�;��*bVm���      �f���H]����0���?�; @O6��^�0�      `2Z�)�ޥ��/zg  �I��k���;      �D�6�{g�M�t}���  zRp�VEΣ2{�       `K*��Trg���f?������ Ћ�;��Z���       &�Zy�ѻt-���Rp�SFVŬw       ���0���7�v�����  zQp�Rk��
       SS�U��3n7���z���� Ѓ�;��*�y�       ��jPpg��^_��w �܁�S�j1�      �>�Ŭ2�^�KW��� �}`�_�      �j�;l�����C��#�s  l��;�o�U)�      Lܪ��1�w�x��  �M��+1���      ��*�2�c�&]�1���  �M��+���       ""���θ��䍿�; �6)��#3��_�      �b��pƫ"����K�s  l��;�7Z�e�s	       �TE�
S��k7�o� `�܁����r       |)wɌݍ���>����w �mQp�D΢Қ      ���������r�ʼ�~�w �mQ�B��{       ^RU�{g�M�v<�;�3  l��;�Z#       xI���4F�ʍ��zg  �w`�U�,�z      �˨"r�;l����;���9  �Aa�y~i      �+�*wˌ�����3  l��;��Z�{G       `��*�-3j�����; �6(�;�2歬U       ��ʡ"g�c��ܼ=[>����� �iJ��N�6��=       ���3��Td\;���� �i
��Nk��      ��Qc�._��w �MSpvVeΣ2{�       `OT9�6����G�S��� �I
��Ϊfz;       ��Έ�o��O����9  6I��MCD���       x8�R��Q�v2���  6I��IU9���      �=S��a��u�d�U�3  l��;���y2      ����p���\~�_^���9  6E��=��a       �ӪZ1�UEƍ��b�  �b+윊�EE��      ���̪4X�Ѻru���  6E��9��E�       �j��Ѻ~<c�  ����!�E�=       �Lpg�N��?v��� �	
��N��yTd�       �ʌ�Y��)'w?�; �&(�;��_�      ��j�;l������  �	
��NiU
�       �ŪwЌ֍��G������� �n
���YTZ�       X����=4�t�e>��g� `�l���az;       �V��3��\?����  �n
��Ψ�4       �U��k'˯� `�܁ݐ��j�;       �R-g���s�&ܺ=_~�7��w �uRpvBU,"�'       �n�Lqg�*"n�m��� �N
��Nh�a       �QU�����w��  �N
�@Y1�z�       `�Z�Hϊ3N׎_�; �:)��U�,�A       R�i��t��l��O<���9  �E��Z-zg       `ܪ�w؄w�<�X�  ��t��!       ��*�M3Z7n�{g  Xw���Ee�N      ��U9�6����W��  �.
�@W-j�;       �`�;curk88��;o� `܁����      `+*J��Qj�q�ڽ�� �
�@?Y��      ؊j9���6����{g  Xw����G87       `[2Z�)����[zg  Xw��*O�      �]�����'�խ�� �܁nZ��       �wՌT��g���w ��Rp���!�      �v����[w��� ࢔K�>*<�      @͝5#u|2���  .J��U:,       ����wF����h�  ��tQ�7       ���Ydd��ng��|��?�; �E(�[W��(       tR��1N�O��; �E(�[W��       ��j���;���; �E(�[W�	       �b0��Q:�1|Y�  ��lUfd�rH       @W�j��;�ۭ����_��սs  ���;�U-r�|       ��2*6F�"�����s  ���;�UU9�       ""��;lF����;{g  8/w`����      ��P1��f��o���; �y)�[��Y�       ���,2�wX��[�kzg  8/w`kZ�<�       �32�b�;����!{��z�  8w`k��C       vJ��%rF����g�3  ���;�5͡        ;�*�e3J�n�� �<܁��Ȩ��       �S��,3�wX����{g  8eS`+�b�       �9�wF���l�ޣZ�� �܁��       ��J��:[e����z�  xX
��V8       `W��X�:�� �a)������a        ;��6��֝�]�3  <,w`�*b��c       �K�ȈTrgtn��B�  K�ظ����        ���m0.��,zg  xX
���y�      �]WU���U�㟺��z�  x
���U�       vZ�A��Q�y���{g  xJ����,*�w
       xECf��ftn�l��; ��Pp6�"��      ���*�3��ݺ�|S�  C�ب�Rp      `/��f�n��Gzg  x
��F�J�       셊�7�s��,�wt�ݽs  <(w`s22�:      �~�V����9`�2���w ��x
lLE��w?       {#�U�������w ���lL5�       �Rpg�N��W��  �܁��J�       �}F���ᵽ3  <(r`c*J�      ���jp��蜞-��=�e�  B�؈�̨��9       �T�ᾛQ��������; ��Pp6�E�E;       {(�"uj�����  ��8�U5�       Σ5wތ����W{g  x
��FT�       ��;oF������  ��8�U5�       Σ�P7�������3  <�q`�*c���       ΣZ�"ý7�r�t���g��9  ^��;�~��       �XF��fdZe|�����9  ^��8�vU1�       .��7�S�����  �j܁�+v       ���o������  ^��8�v�w       ���o�������  ^��;�nU�       �ZU��s�:���� ��(��9��      `�UdD��0*��f��#���f��Uy�      ���(w����U�̓[�w �W���U5�       �C�n���V��; �+�	֪Һ      �X���;��{g  x%6��ZU��      `ZyŜ�9=����  �JQ���̌��       ֢23�=8�r�t��  ^��;�6-�/�      S��;w��  ^��;�6�|�      06�_è�ޛ͎���5 ��lT�u��       0*�����_E�˫��; �˱֦�)       �M5��3:�9�۽3  �eT`m�k
       ���w�������  ^�8��1DE��       kU���>�Q9=����  �r܁u��       0J�܉3.wNo� ���|��I6       F�f��:ݹ����  �rR���Pp      `�Lpgd���h �Y6��Z��y       F���N�Q9[e>��կ� ��|k��      �XU�;qFg���� ��|���c      ���� ������  ^�B*pa�Mo�-      �HUd��㲺7G�  /��X�T      `�*RφQ9��zs�  /��������        Uz6�˝���{g  x)6����`�;       �VQz6������w ��b�\X��:       #W5�gTN�Ƣw ��b�\��;       �usF���l8��z�w �SJ��G<       �f�cSq��ɻ{�  x1o�B*c�Rp      `�*2��8�r�t��3  ���;pQ�       &"ݑ3*g�ûzg  x1�n�b<�      �D�;rF����; ���tRU�       &�9cs�4��; ���t��;       l����Q9;� ��܁)�       ᎜��w6,{g  x1�n�B��:      ��pGΨ��a�; ��)���      �I�ҵa\���M ;�8���Rp      `"��#wO�h�o���굯� ��܁󫴆       05����?|[�  /d��[EYC       ���4��Q�sZ��; �)��Ve      `b�08ƥ���; ��p�~�      ��T��θ������  �B
�����;       ���θ���7��  �B
���U>�      ��֚��rwU�� ��l���Pp      `Z�]9�rvox�w �Rpί�!       LK����{gòw �RN�+��G;       �R�oè��r�; ��p�R^]      `r22Ӆ9����:d �N�9�%��:       ��LqgD�V�����^�; ��l�뙻    IDAT��s�2�      ��2���9���zg  x��;pN~�      �D
��ܽw��zg  x��*p.&�      0UU��12��;{G  x��6p>��      �D�3gd���-�3  <O�8�      �*��{�ۛ{g  x��6p.��;       S�ΜQY��/� �y
��y�X      `�����Z��{g  x��6p.U
�       LS�tgΨ���5�3  <O�8/�       L�;sFe����  ����O��u       �ɫ����8� �y
��C���ct       �+#������E�  �SpZ���       L��s���j���  �<w��U�H      `��n��5�� v��	��*�
      ���pw�h���G ��ᕏt       ��X�A �
��y�����]��Xr��fVUw�
���ݟ�6`�B�tU~�'|1+Y�������C>��� ��)�      �o��1��E���u�= @����rH      `�*ʳs��O��{ ��;�)�       �G�����  w�S�      ع����>����  w�3J�      ��yt�X���= @���gt       v.=;g0-_�k�  "��'TL��       웯�3�yi��{ ��;        �N��p�{O  !p>�1      �}+���r���{ ��;        ܬ)�L��S�  "��'T��      ��U��j�; �
w���      �ΥG�e��k�  "�        p;�L[B� ����o�      �s���e�z�= @����rH      `�<:g,G- �
nJ�[M�        cYZ;��  B��h��       �Ѥ� X7%�M��v       ��,Z2 `ܔ 79�P�      @Dd���*�% ����I�r�=        ��Ti� �UpS�$��       Q��;�4! �*�       �3���di��#  D܁M���       `0�^�  �A�        �w-� �*܁�x[       `<KhB �u��Y�       z`F�5iB �UpS��p8�       �;��� �w�&��       ���(M �
�� �b�;0���m�=�Y�G    آ��?\{�@_Ǘ���3 �[F���� �J܁�,�� �'�c_��    �?-��?Y6�@*+���#]� �JU����4         �c܁�,K�       0���= @D܁Uơ�       П�3�tM +!pnҖ��       �W�2l� ���7yy��       ~Yvm�5  ܛ���e�*�       2lp ���79��       �_��� X�*p��W�W       �" X	�;p�i�       Qi�5CqA +!Tn2����       �]���  �O��d��K�       ��� �#܁�,���       П���xg X�;p���kD�       �jQr`  x �;p�6�^�      `��  A�ܬ�!      ���  B�ܬz        �yx�h�E ����YFx       ` Y
w `���J�      ���g�� �����       ;W��9  <���Yk�       �[U�	���  �J܁�y      ��+��  �!��g8�      �s�3��] `��ͼ�      ��U�g�EH ����f�       �[��h\� �J܁���      ��5�� �!���*�      ط���}M� �A�ܬJ�      ��5-0CqA �!pnV�o       �UUSX�P\� �z�T���r�      `�2� ���7�&p      `�*b
�;CqA �!pn�|f      �����D	 ������       �\��p  �w�f��      ��i;CQ�  +"pnV��>�      �N�  F�|JsX      `��3s  x�;�9�       ��� �������      �N-M  �"P>��a      �}�̜Ѹ����R��g       �ZɁ� X�;�)�x      �}Z���  D�|J��.       ;U�v  x�;�)���      �UMM�  #p>ei��{       x�V9E���+�E �������|       �CYS�  E�
|Jk�{k       �N���#s�� `]����K�       {��6�� �ڸ�>)��q       ؛��� �	܁O�H�!       �J�ep� ��8����o       ��xV  ���Vu�=       <S����������V-�q       ؕe���������k       �IEekj`�� �F�
|�R�7      �����z  c���f/�      ������5 �����y��!      �ݨ��.8�.i `e������      ؍V�3����?���g       �g���  ����~Hk�w      �]X�c�I `��t?�y;      ��hM�`\� �
	S��Zz�        ϰ��34 �Fw��4�w       ��jZ�� �����[�      `x-�P���{�� �B�T��,sL��       �����8�ѷ k$p~�<G:�       0�V:F� `}�x?&3�o	       �k�g��VC `��x?��8��       �5���� X'7��kUw       �6���`,o �ʍ7�Ö�~K       Z[���% ��(�a�6�      0��8�R3W4 �Vw��->�      ��ZձU�)��� �J�R�v�33�Q      �1�Ɔ�����r��AF��{      �����3  �^R���J�y       ��,FS�Y��  �Un���hK{�        �0�N�  �7���b^�w       �SQ�,b`�b{; �fw�.��~O       NU�  �F�
��u�)      ��Tš�w�� �L��Ų��       �iKz�   {"p�ɡ      ��,��a<� k�����       �eYR_À��   ��8p7�R��3       �=]�v]3��� X5�;p7�9mp      `�űYt  O%p�f�s��+       �PQ�*����� ��	܁����t�      `m)_2g8� `���]�J�{       �0Wjk�� X97��]-���g       �{Xfm�ѷ k�&��y	�      �<���d��  �w	܁��      0�V�Қ��є� ��	܁��\�Y^�      `Ӫ���oF� �܁�����m      `�%}�  :�wWK{�        ?b^J��p,p �@���"p      `㮳���� � 7���]��      �Y��qn�  ���8pw�u�"�z�       �QGO�Q� X?�;pw�U>j      �&���g�{�� �
�;��ű�       ��w�cU! �w�!Z	�      ئyI)0�qQ [!p�|-�;       �SU��U��x\� �V܁���y���=       ܢ*�v @?w�!�e�,_�      `[��b9C��� �w�a��       lʼ��po�v `;���,K���       n1�z��  ��ܐsY&o�      ���q^����U l��x��9���W       lBEK
̀�e l��x�VY�H       lò�/�3(�	�����z�=       ��Y�Θ�' �D�<�u�      �~��뤥a8i{; �1nʁ��\��3W       �]U[�=<��� ��܁��\s�*0       k�,���$p 6F�<XFk�        �ڼ��  ��x�e�c�       ��\���aH��{ ���1�rM�;       ��Z�sd�9��2�� ��܁��\���       �kZ�1���e l��x�VUu�=       ��6�g�)� �	܁��/�g       �_s���{x}; �Ew�)��;       �SU��2�Rf� �fw�).�<F�S       �Ҫ^=�fD�l `���S�Kf�/_      �.˜��3�C�4 ���O3�x�=       �G�9��g�GH�; �Qw�i��z�=       ����.�I̐\� �V	܁�9_�Y�{       ��h/�b3�L7 �Mw�i��[�       �ǲԱ���v `���S�%^{�        �9�)�  6L�<��Rw       ����r�3&W6 �ew�.����       �[�z�R3��=  ��	܁���̨�      ���9��g��(��M�O����{       ��2����v `���ӝ���SX       �RU��%d�Ʌ l��x��%^�)��s       �O�ŋ�Q�� l��x�VS�V��s       �O�Y3���= ��]\�z�=       �t�ơ���v `w���5_"é
      ��j��5���.l `w���9Y�z�      ��,K{�=<�W7 �܁N2Z�?       �T�k{� �S�  �aw����z�       �~TD�.��aHe�; 07�@7�s�L��       �Ck�Z� fP.m `w��y����      ����3��Lw `�R���Ro�g       `.W�;���� �>�;����/�NX       <VU.W;�W���A܁�.�<f��{       ƶ,���(�v `$w������?"       �P�9^z� �"p F"p�;]�-�z�      ��*O�I'ðRw č;���<�LS.��       `L�R�UV\3��� ���n^2�V��s       0��/�g�G� ���p��[�       �霖�1,}; 0�;�
�K�FV�=       ci�^�&f\��{ ����p���#       �ni��{x���� 0A)���,��{       �r:��� ��X��9�"�w�       ����:I��� ��X��9�SF�=       c��z�=<�=� �x���d�s���      �1�/��{x����� ��X��%޼]      �L�Kjc�� ��x`UN�|�2Z�9       ضyno֫1�I� J��JE���'�       �!�kz���2�� �I����oa       |VM�K�b�� �y`uN�xͩ��s       �M��U�{xW7 02�;�:���ŧ�       ���5<sfh�p &pV��_"���       �IE�锇�s�#eJ* �q	܁U:��u�Xz�      �����UXo͸�� ����*��bY�[�9       ؖ�5_z� �4y ��X��ez��      ��d�震�c�C�� N����)^3���      �mX�z��ޚqeV����	܁ժ�X�z�=       �p��k����� �܁U;_�Kd��       �����9�0-� ���V��4#J�      ��j-^�~k�V�)�  �'pV.cY��       �����g�G�� ��;�z��^A      ��UM�S�`�$p v=�z�sB�      �o��x�ޚ�ej' �}��1_�K�)       X��%^{� �$n �D�l��%_#�i      ��Ҫ���d};C� `O��&\.ӡ�       �ϲ������ ��܁͘����       ���)_z� ��Q��� �~܁�x�ȷ�b�=       �PU/�9-�fl�p `g��f\�i�*�[       DD��Ro�g�G�� ��E�M9�۷��      ػ�ʏ�t�=<Z�N ��;�)���u�r�=       }�%^[Ym���� �	܁MYZ�4��      ع�%<;fx�w8 ����qʯ��e      ������<�^�� ���6�t�cD8�      ��u����eVX� ��ؠ�뵾��      �>>N��{x�I� ��ؤ����S,��       �Z��<����Ud��= �Ow`��˔�ձ�       <��o�g�G�
 �gw`�N��^W      ؉��N�<��M� ��ج�S�N��       <�2�[��ѕ} ��	܁ͪʸ���       <��9^{� ��i�; �ow`��?�W[�      �ת^.�I���\� ��	܁M�\S��[      0���z� ϐY�G  �J
l��R_#�       ����Oy�=<ZfEZ� ��ؼ�iz���{�      �c,s���7{ n �XZ��      ��>���{x��L_� �C��_s���       �WUΗI����/�  ���?0��e:���      �r�/�g�gH� @D܁����-2|�      `��|�=<�� �w`�?���Xz�      �},s}i��ǀ�ˬH�: @D܁�Te�s}�=       �P�q�^{O� n ����P�ķ�lq      غV�z�e��Ô�{ ���C��S��^z�      ��9��K��R� �W��p�O�-���       ����q�t-���;  �A ��<{�       ��]��%B����  ���P��\�"       6'+�L/�ǀgH�q  ��;0����m�r�=       ���xk��e&�: ���Cj�q��K�9       ��霯�g����uz ��L�����Y��       �1���|I=�`{; ��s  �u]��*��       ��9_���,)p �Uw`h�-�|�      `���S{�Q�)g  �5w`h�|���{       ~��ھTYi�>L.u ��$p�q>��"�k�       +��1����%' �o��{��ަ���       ��y���Yi�>dV�� ~����2�����      �P��G|�=<ˤn �]w`~~�oӔ��      �̲��u����� ��;��2�<�[�9       �k��,��� �}w`7���O9��{       ~Ѫ^��I��n�V ��� ��e������s       ���S}�=<KF�� �܁]�~��"���      `�Z��t>hW؍�� �qH v�|>���      �v�ė�3�3�~{{�� �B�	����~�,�2      �~��y�=<Kf�~��t��{ ��;�C��e�gF      ��].�k�'��Ǵ�˽� ���ء��S|��i-      �g����1�����"s��BN ��;�K�|�(3      �'����j��>6��=""���   B��TU��Z��      <QF���x�=<���GD�o �A�����ӗ)��      ��\[}Y�\��Ȭȍlpϲ� X'`�Ze\.�5,q      x�����|�=<Ӵ��=""C� ���ص����4]{�      0����u��.k����,�+����6/�׹}qF      x������{
x�iCq{DĔ�	 `Ц=W    IDAT�������SN5��      `T����:veK��#"b���  w���)�yz��      �*�L���+�����͔i9  �
w�������)mq      ���՛���ʹ��="b��w ` �-��9���      pO��[�)�*2��L���{ ��;����=~�&��      ��e�������������{ ��;����)�ײ�      �.*�O���79m�;�,��U��?��-�       w`{;{����1e��Up� ��%�zm_mq      ��g��ٟi�u{D�νg  �����ߧo���      |����r���}ɨ���B�i
�; �
 �ɼd�s��      �)�i{;���W:2��  w�_��{|˩��s       l����r�z���6��="�ө�  w�_5/S�s~��      �����l��=""s���3  D�~�����4��{      ���e{����g�������!�o�  "� �i^2�װ�      �Ȩx�H��ٝ̊ൎ���z�  !p�]?��O9�-�       Ǽ���:B������= @���w�e���Hk�      ~[�������ɨ�#)����{ ��;�������a�;      �o���r�G�c�H�,8O���  w��kY2?.����      �odT|�>�����"�AR��"���g�1  "� ����kdk��       X��5��m�=���L1ʅ̪?�9}� X�;�P�����;      �_TT��{���.e��="��? l�����1�E8�      ���U�����̊��[�w `E� X��{��-�       1��^z�W1�GD�� �j�n�q>�D5��      ��}�뛕��Q�/�Gr|���  �F���c��~,K������Ǚ��9�9MK��#��[�F�/ �e)��Id[�8b�"����(p��Nفɶ�ȑPR�'E�lQ�������}X_.�C6��3}��o~?�7�~f��Zk}�z�&��%�s       �Rk�ONJ�uh��a�j�_�Zg  x�^n\�����g�      ��ur;�3@u���#"�M[g  x��;�8��R��      ���u��d�����rM����y�: �{����b��Yf�n�~oe      <\��I�Nm�(k���/w `i(�<��q�w      `�,�5���5|���\�~?�Zg  x��'4_dNϺ�H3�      �&�1���v6T�Rַ���;�3  �G��)Mr;3�s       \���n�����p��70��o� �=
� O���g�^dt��       \�G��j�Z)�����^��Zg  x��;�S�˨��;      ������U56Sf]���u��: �{�y <�Ǔz%K,Zg      8o��r4.��9���������X�F�  �Qp8'ge�u]?b�?I      l�����_x�{����t��u ��(����㲟��[�       8/]���i��:��	��^�w޹���9  ޣ�pNf�,�ilG�q      �A��8vZ��V26c��7�]�  �Sp8G�㲛��9       ��|^���Mد�+Ҭ��u�V ,���]͘�t����f      `eըy8.[�s@+����1.f�3  �O���MN�VD�b       ����ܩ�=�`���� OZg  ���;���8�A�X�N      �j��x��9���Yo�����  ��pΦ���wÈ͹�      �A��Iݍܠ�jx�ކ5��ø�: ��6�r����^����      ���:�}6�f��GD��_��  p?7$ d��<;��"͸      ���x���)��M|��?��m� �~xIpy��eT�*�      Ko:�۳Ef��N��a������[g  ���;���q<��,�h�      �j-��2lZ*��zG�_n �~
� ���E׏ؼ��     �UPc|�56��5Jټs�̌���Z�  ���;�%8�A��u      ���蟞�^��R��հ�u���i�  ���K3��5��<�v;�u�^�      �X��I�Nm�(����[�:o� ���.����E�       ��c{6/�:������Aw�: ��m����5�xR�d��     ��j���8�Z瀶6w�="b8�&�3  ���;�%:9+�n��ͽ9      �ˌ:9����l�M^o����/��  �~~�p��e?��[�       6�lލN�J�uhk���#"�[��Zg  x?w�K6_d�Mc�dt��       ��f��qn���0�����k� ���8�F],�*      ���4v����F)������o��  �~�V 9:.WJ�y�      ����Oʠuh��5;[�wZg  x?�j �Lg��fu;2�      \���� ���tT��e����˭s  ���;@Cw�s�dt�s       �o>���y��9�5���l�E�  �r��Z3���A(�      ��s�uh�z�{�[���  D�����ޠ[,n�     ��Pc<�{�o��ߴ=�ƭ3  <�K6�%p4��eT��      �ݢ���i�a�eZo���V���  ����/2Og�]�,      ���Q��8�[�eP|��[l��i� �A����"|      8/5���΢S��߮�U�Q�  �`idǕRb�:	      ������'�A��������K�3  <��;���J���Nd��8      ��2j��n����?@����ϴ� � 
� K��8wK֮u      `u�����"mVCXo��V׽�έ��� � 
� K�֌��y�Wb�:      �zj���Z�e`����F��u ��QpXB�i���Nf��      ��q��v��E���vF�q�  �����s72��9      ��q6�vg���Q2����[���  �0
� K�֌ãz�����      ,������2h��E)��f8���u ��QpXb�Y)�Yݎw�      �:箹j���c��3�_n� �a����q�     ��:�՝٢h�CDDT��bk�k�  ����j͸{W�ļu      `�t����9l��EO#�zY��Xp ���9�0��2��vdx�      ��q�Fo�������?�h����  �A�V�ݣ�-��      |�t;�y�n����Q��>��p~�: �qI�"j͸{\���-Zg      ��j�?ǰuX�a��l�����  �A�V�tV�l����      6Z���Fo�������٩��u ����b��n��Z�       �9�֝�,�y��JV��hԯ��: �QpX1�f�=��z��Y      ��Wk�OʰuX&����v���  >��;�
��J9�u��a�      6HF���؋0��)���<���?��׿�: �QpXQw��ND�{�      �_����;[U^���z�#���N[g  �0
� ++��(�����I      ���u1���s�2�i?=����u ��`���Y&��A�X��      \��w�b�u
X&5�z�c���~�u �����Ɠ��bQ���      �Pf��I�몚|S��G�m��WZg  �0.� ���qdZq     �u4���ӳ^�uX&�a��	lf�u �������q���Sr     �5R���uX.5�r�cˌ������� �a����Y��g�Y��     �Z�q<.�5�uX*%y<��������I�  F�`��=ν��u      ��M��t���-j�b��I��,�Zg  xn� �H��G�J)ݢu      ��u��'�A��lz�NOlw7~�u �G�`��楜��nd��:      ���Gǹ�:,������h���  �(����q�j%=      ����؛/2['�eS�T<�+����: ��PpXG�qx���u      ����utrZz�s��)�۟J�5����[�  x
� kj��O�,ݢu      ��Z�e�:,��(�?���b��;F� �ՠ���&�e���03��     �R�q<��Z�uX:=�������: ��r�����~dXq     ��U�lZw�fE��'�F�M������v�  �ʍ���5��^����      ,�����7l����>��h��?Zg  xT.6�t^��I�g��      ˥杣�m��Q����2����  ��;�����żFVw�      �2��$�kU߀����akP����~�u �G�	`cd�9*���k�      ��N��ٴ�n���s��;��  �8�$l�Z3��,1o�      6Y���Ѹ[�e�Y����y�߯��u �ǡ��af�RNN�~Xr     �V��Q�˪d��e��J�  �C�`�'ek1�����;      \����U�x��5�z��:����3  <wK ��Q��v      �Tg��9�}x��8�>O�^���]���s  <7L �F��Q^���Y      `t]�˰uXN5z�L�nwgq��;�  ��� l6�rr�DF�:      �����8v[ǀe��i����.~�u �ǥ����'��b^���I      \���uoѩi�Ô���"����h� �q�s ��^D��       .��,v�f=x�Rjd�kjwX�F�  ��� Q#��(����Y      `�t���e�:,��%�]�~/j�O\��Z�  x\
� DD�l�e|�d��37�؏      ���5��n��̊�����8}�vN[�  x\.���Io������C��ܧˠu      X]5��s�V�x��5�z���r0���  ���( ���v�_ً�������      ����Y�Ng��U��������j�  O ���%&�9*�w~��_x�C7      x�E�O|1>H�I�~����3  <	�� |õ+�?��"''1�Z��t�v3[g     �UPk��=*��9`�e�ȴ�~���_�S��z�  OB��ox���FFD�Y��:�������p��q     �R���q�E8[�R��/���l�: ��Rp ""vF�[��ӳҟϻ�����&�v�     �aj�'�?_8U�RJ?%��n�;�3  <)w ""���22�}J��4�5^��ۯg�E6      Xn5N�b�lZ�0�dV��d{w�3  <)7V D���+~E�F�d����~��_z!{�      ��|QG�2h���r�%�;��_�� ����>�1|�z�{]��$F�����,�+>      5j��Z�eWJ'͗cgk���/]���s  <)w������a��2�Ű?���*í���      �	j�<<ʽ��>PF��~���M�m� �i(�l������y�'n�g��({�����2�v=      �*��xR���f�aJQn�L������  �4�6��7�y�d[��|�f�>};      �X����{6��]��(���@.�����[g  xn� 6��k�\��%��89ɭ�ѽ�J�_%��      ��|^G㓞1(�5JZo�L�^��?v�?o� �i(�l�O��d��/���I�JD��ۥ���s4      XJ5j��Z�UP4�.�������9m� �i���P{;/������"�t^����ϔ��+~�      ��j�<<ʽ�xI��TJ���~�v�o��  �6�[odD<ݓ�ӳ�_,jo0�����pgۓ<      �U��8��t&"�FQnob�`�3  <-w�4D����y�69���"��3��2��=�     `�dF=9�{g�Գ�GP7����u ����`���~�|��kdLNs�Q�Ճ(���ڬ      `}ԘN���I��:	��Rj���&v��/����: ��Rp�0�D|���m�/���Il����g���rp�       4�uux8�m��� �FQno�ڕ�W[g  8
� �c����z�����Y�JD��ǳ��+i�     ��Vk��Q�iVE�Dj��A�B�  ��e%������wۿa>�2�ǰdv��]�/ފޅ�a      p�j�=νZ/�|�I)5�z{;Yb0����1  ΃�;���LƵ+��~�ӳ���_J��?SW��]     �jɈ8��|����2j���vG��O}��Ϸ� p�6ȧ޼��o���9d|�se��}��z      8?5Ƨu:K�
xD�(��v�`���3  �7c ��Aċ�]֟�1��(��Q�>W����;      �o:�����k�VE)5|렽+���: �yQp��_/Q��-�ך19�QfԫQ�����     `�-u�h\��s��ȬQ�z�2����Y�  �E�`��">������.��$�Jf�̍�}�39��>      ˨��ݣ�n�V�r���u�/��՟i� �(�l�O��Q�孷�o��rzV�Jf�����O�E      x�Z��qٽ�"���g�����k�3  �'w�5��E��Jۧ
�Y�f�:Ȍ��W����o      ��F��q�/:M]xT�5�z�Ҹr��j�  �I�`ͽ�r�ְ����i�E�̬��d��R�Zg     `�՘���l^������+������쯴�  p���Xf�[�/˳���ilE���]�Q�=�~     �FF==���g�0<��Sޥ�7���|����u ���`���\��^����Ԛ1��(��,5��gsx���E      \��i������*)Y#�z�2�vu�{�3  �7�B�5��7����]9��v�����/~�ww���     ���/���l����F)��������Zg  8o
� k��Ոgo,gq|�eNN��G����|˙     ���uѿ{T�[�U��2Z:����O�� p�\z��O����?_dNNcT2���(_|�{�֩      Xg��ޝ���K�XJ�ȴ޾l�w�g��n�Z�  �m�ۏ <��툏��:Ň�ϳ��խ��]���p�g�      \�Z�rx�{�:��ǑQ���et����[g  �
� k��32Wcvb:+��2��x+zo���     8O5j�s�p�K�}yl����  .��;��"^��j=�;=��b�̬/$�����     ���c6/�u�K�Wjx-d9�zYw�?�: �EPpX3���1��z��&�1�Z2�~�����     �j˨1>��g����d�L������l��;���: �Ep�F2#>���]��$�j�2"�;?Q��~4{�S     ��j�Ls���8s��V#�r�2�vu���3  \w�5��3vwVo��=�f�'9ʌY��^~A�     ��7�՝�$�s�*�X݃�qp���[g  �(
� k������֌��K�5��L��\�}     �#�/��Ѹ7l�VQ)52��/�Ѱ��ҏ]�+�s  \�A�5��͌���%�Eyr���e��=�-Ûו�     �p]Ww�r�uXE�5�r�һqe��[g  �Hʂ k��k�m���"srz�������w��� ��     ��Uk��Q��z�B�%�Q�r�*�z����  .��;��ߍ�ȭ�)��|����n��n8�������      <@�ʻG�_��$x��ՐU���;����s  \$w�5�ֽ���|�0���tV�%��ގ���#�    IDAT�.���z��     �j����s�O�d�L���`ov����WZ�  �H
� +nk����������g�:Ȍ���{?_���z�3     �hj�<<���< �ȬQ�r���yu��Zg  �h
� +��W3z��_4?9��b�̨׮D��۹�Wr     �p5�ǹ?�G������rp��w�3  \4w���E|���nr�n%3�kQ��w��7     ���q|���Y:1�'�+5|�`u�QG���: �Es���^y)c�����ߔ1>���FfF}�f����e�     �fɨ1>��gg�k�VU�i�}�ܼ:��;�s�: �ESpXao������8F���������2Pr     ��Q'��wz�Sn�'�Q���Us���g[g  �
� +���2�l�z�7�{K��u�����w*�     ����uorZ����*Sn_=W�ϵ� p�V��76��]k��$G�Q#">�R�?};�s     pQj�����Iq&O�Wj[=׮��_��W~�u �ˠ����D<�l��՚1��(뽒��d�So��     �54����7l�VY����Wэ���  pY�V��7J�ީ������~s����9�īJ�      �d��F��e�uXe5JQn_U7��u �ˢ��b�G���:�rYt��I|�����,��>��ֹ      xz��ۺ{XF�s��Sn_]{�����?�� pY�V�'^�(i���]��$F%�����?U}Q�     `�u]�=,ۑ���i�J�c��1���  .��;�
��"�����XdNNb�dt�5?��2xY�     `%u]��9��j�	�J����W����W[g  �L
� +䵏e��}����K�q��������[��     �Bj�zw�r�VGc�42j��ܾʆ�����_j� �2)���̈�^� �Q�YN��U"�,5����/<�~�     ����a�+���Rn_�\���;�s�: �eR�X/=���c��QMg�;��V�{%���l>���;     �2���{T��X�V��Rc�ݸ��[�3  \6w� +���<<��,{�g���{��_��2|憒;     �2�Q{ws�����*Y#�z����>�ܕk� ಹ+X7�e<s�z���ɽ׫����፫~�     ,�r�0�-���ˬQ�r�:�~����w�Z�  �l�V����m�Xr�����/�]�ו�     �B�Z��~�9��W��ܾ6n^�?�: @�} Kno'��Z�X}�J�u�dt�A�?_�W�SR     ��j���0��s8=M��Q�����G[�  h�e-�������9���7J��a�};���]     �B��+��y�����ō���w~���: @J} Kl0�x�c�睧{%��*���V���]�J�      ��r�B��CI��us����Zg  hE�`����~�z�y����K��,�_9��     �2�Z�]�v87�5JQn_'όꏷ� Њ�;��*%⓯z�wQ�_r��o疒;     ����F�ܾv�]���ܗ��_�s  �����>��������4�eo:�C%w     ��P�ݱr;��^���~���Pn 6��;����k�B\�ӳ쟞u��     .RF�=����9���R#����̌����m� �%w�%t뙌W��_��|}�=��     �[F�=���p~J�r���v0�ԗ��|�  -)�,��ox�w�Nϲ?��В;     ���Q��a=�ϋs8'�5JQn_W�^��r�  �)�,�+���:�f�Wr��     p.2��8��v8?5z��k+kč�c�s  ����d�z�D��!_#�g�?;�[�/���*�     <�Z���8�ϝ�������Yk7�-��O_�?[�  h�e/�mE��R���J�������F�u&     �UQk-w�s�Pn���+�����37���: �2PpX"o��Q���e0�e��n���u     �UQk��9��v8_%�r��ˈ��>���9  ���;����">�q����l���i���     >\���9���s��)�F)��������_��[��: �2PpX����5�޾l��,J�      ��j�ݻ��U�]p�j���7�s7��k� `Y(�,�̈�^��oY��Y&'J�      �u��(��r;���f�F���^�Z�u �e�2`	��\�����e6_d���v�Tr     �����v��R#�z�&�q��Η��?m� `Y(�,��ox�
���ng��H     ��[tu��a�*���+�ܾIn^����  ���;@c׮D�z�u
բ˜Lbd�     �d]W�ws'|��]f�R��7Š���Z�  X&
� �}���z�J�%w     `s�u�ݻ��p2j���7ʳ7f����;�s  ,w��v�#>�b�<�{K�9Rr     6G�������H�v8��7ѭ����u �e����'_��4m��]�X�     �5f��=*��I`]�JxwdÌFu1<���s  ,w�F��7^�tb�u���3S�     X;�Q���sx���Wj8n�</ܜ��w��y�  �F����>�1�[o_]y<��Zk*�     k%���v{G�ްuXWE�}c=s��[g  XF
� dF���n�:�5�x�nQKfx�     ���'u|��N�*�FQn�H����#W���9  ���;@}1cw�z������b=%w     `��8>���i�N�*�F�8V�T�ݘ}�u �e������u��W��4��Y�̮u     �ǖ5������ZG���ܾ�JԸv����9  ���;�%{�Fƍk�����Y�O�u��     ���yxX��O F�}�ݸ1;��/]���s  ,+7� ������t��ӳ���     ��Z���<�-z���JD�)�h�߬�u �e��p��w#^z�u
.�t���i)�     ˬ�j���<�/�n���[nϴ޾�������O�� ���.�[���=�0�y��I��O�     ���uup�(���.R�Pn'��9������� ���.��0ⵗ=�T�E��$,�     Ke���=�ݪ�*�F)��D<�l�OZg  Xv
� �䍏g�z��7�b�9��%w     `	Ԙ/�ѝ�޶��ʬ�Sn'"v�?��W���9  ���;�%�<� "]��8�[�      6WfԳYݹ{����N���ݺ1���  V��;�%�����W�q�䂨5c<�Q�jf��     ��ɨ'�u�x����FQn��J�8�?���9  V��;�%��_��뿩���K�'��-j�'     ��QcrR�'e�:�����c�4��1��~��/�� �
�.ٯ�Z��/�܉�����|^�%�k�     X_5�<���i������vs�>�?3��[g  X
� ��ֈ_���䷬v�qrZ�i�%w     ��ըyxg��# N��o�=���֕l� `U�yh�ֈ_��.~�w�ܹ�t�����Pr     �O��w�0���l�6AI�v�ݭ�g���9m� `U(�4Rk���r��ܹg6�2>�mK�     �ӫ�uu�w�~���e(Y�ǿ|�̌oƏ�� �J�꺈���]��W�ܹg��Ob;��	     �I՘�c���܍Pn�ː��<�����/��՟i� `�(�����,}κ.�g���~M��{]��8��F��     ����4v��Q�r;\��=�v����u �U��<�~��}�s7_D����������=�fOb��w=k�     ��Ȩ1>���[g��Q��s�ǃ��]��3'�^�  �F�xl��0*}�f��������efޓ19-�٬J�z     �p5k������Zg��a����ͳ����¤u �U��<�������"���+��N�J���n)�     R#��aLg� ��W"2[�`iՈ[���l�  ���-��J��z��Nɝ�β79�#%w     �~]W�w���|�f��(�����;?t�� ��܁'�q��z��Nɝ�/��O�vz�     ��Ţ�z�0�����I��G�³��n� `U)�O%��ͻ���{���w������$GQ#�S3     �H�Qg�n��Qo��,pY��y�Q]���W���9  V��;����[�XO�Y�����;�j�E�'1��Xs����{��������׾��.�. 6��؉��I���t�&�N�zʤ�'61&�Ǯ&Ů=�4MۙLo/2�d:���M-c@HB�27�� ���{��Z����`�$Α��Ͼ|>3/��u�}�����   8f2j<�Nn�}G��)�s�n�~�ѻ�+��� pX���"�,��K�<����8V��̮�<     �~�����x��w8nZV4�v.Cˊ����� �0Spv�Nɽ�G�t[ɝ��1���tڭ�%w     8ª�vi3�L�9�;7�������p����g�; �a��
�*����v�;����M%w��t��q�Yr    ����Z���N�-����7�f�����S�  ;w`�5%�=3�F��]J�|��"�p�YQ�ލ     GBF��څKy�+�v�o��\��'�ۿ��s�m�9  ;w`O��h:�{b2����x⢒;�l�En�b�[T��|     ��V1w'/m�"��a�e(�s�n�n�`�  �w`ϴVaHzoL�#��`O\Pb�UdǱ:��R����     \����a�N�}g��(�b0p˕Y^������� �(Pp��@�}�l�"���.Wr�[d�'�<�֪�;     :��f��Κ�|�AFE��γp�u������B�9  ��{N�}�l�"��`_~\ɝo�=��h\�J�     p8tK�/����e�Y�x�'�T�w�̌[o�7�� �Pp�ŠU�����#�}O�}�̷�/2��X��H�4    �)3j����d�f-��b�B��g庳�K��3�~��  G��;�o%��2_D���.���o��"��\���!     0�I���lk��П�r��4�������}g  8J܁}�ZE����"⾇�xTɝ�P�1��|V�-��;     QQ�5���q[�;g�V��<k�����~S�9  �w`_e�,�+�����.>�E0Om<mK�i�*�    @ߪml��鬹��)��\�r��3  5~Q�]��!����躈���g��Զg9�k�e(�    ���Xt�|�b��/2�NǙr;���RW7_7���s  5
�@/2#��3U�~��ONɝ�6_dn�r=""�s     �"���:qq�]U���)�vv�-7l����W�� pԨ���,K�{�*����.0O��"���6��R˴�     {l8��[��J�9�k��<g-*�����s  E
�@�vJ�}�8��"��#���;O'c<��ɴV[��;     쁪j�6��d�}g�㭢eEk�Oy�w������;�� p������>�ɊG>R��C�m�r0Ǻ%w     �M]W+6��|Ѳ�4pܵ�vvͭ7�~��  G��;p |c��a�^�ħ+�`��;Og���։�*='     �e�t�N\�h'�tۡo���MלY������  G��;p`|���^���T���U��<����8Wg�Z��     �V��V��V�N(���n�~����  p����N����^���+�{��Sr�ieL�mi4�����     W���6��t�������첫Nt��s���  G�_��G�}�=�X�;�]1_(�����l�Q�gFe�g     �IF��z�R��/2���{fo�v��;�;�}�  8�܁�A��{�o{W��Lɝ���2��b�[T���     �Sɨ�L�䥭����;g���ru��r���� �Sp,{��o{W�m�e�^E�p���Y,����<     p�Tn��pܖ�N�p��^����G���y��  G��;p�9x�{�/E�s_�C%w��d�K�I��L%w     ���j��f�ޞ��w8 �1�W�Qg���  ǁ_��/��9��S�È�>���%w��|�m8�������     p<e�l^k�7��b��w`�r;{��'���7��s  
���Д���x�Sr��J�<�E9��b^k�     ?�q���jk��pP(���ZT�pM��s  
�������go{w����;Ϭ"c4ɕɴV[��;     �BU���83����� ߠ��^��y���7����s  
����������ŧ>��η�=��p�Q��    �hʨE׭\���g�f��v�\E�r���c  '
�������"�`�d����]��V�/�5h���    8R2*��:uqcp�B��v���޾��v�_�� �8Qp%%��W�W<�Lk�<����$W&�ZmJ�     U��V�M�R�Q�o���~����o�� �Qp-%���OW<�HE��;���,�q�gFe�g    ��)�]����ӳy3��r;���3������  Ǎ�;p�)��������:%w��E����E��    p�dT��u��F;Q���r;����G�  �#w��Sr��>V��*��
�|{�q�L���"���     �e�j����hҖ��|+�v�ә��������� �8Rp�%������{��bs����ٞ�`8��̨���     p0eԢ�����l�̶����~������w ��J�82��}�����8Iɝ˳Xdnm��b�2=7     ,��I����NT��A���~�j�fW�N���  Ǖ�;p��ח�n��d����/���<�I[�Nc�et}�    �'��<=�r�A����Nn�y�����y�9  �+w���Yr�;��7�G��]�韕�$.��,�q�gFe�g    ��T,�Z9)����f	(o�뫋ŋ���}�  8���I���Î�T��+>�q%w.�b��5��nQ-�)     �+�b<��.n�U�w�i�������l�����4�; �q��Yi�}�|���@U��2��*c8���i�����<     U�.mřѤ-��x:;�v�v���V��OL�N�9  �;�O�HK���7��lŽﭘ/�ܹ|�YG�Qa�    �=�Q�y�v�R��͛�v8�Z�Yo�>�y��7��a�9  �;w��Sr�?_�r���U1�VT��-�̭a��f��2��    ��2+��8uik���Yk��No�׺�����  (�Ǆ���y�B�=�w����ΕȘL��h\k-C�    �]P�u�t�R��Lr��4�3(�ӳ��4}ϛ�t�f�9  Pp�%����q��]|�q%w��|�ms'�����     �,���v����Nλ4�\k��N�V�����3��  �Pp��o�����v�����g>����Teǹ:�Ɗ5w     �TU�66��p4X�;��Yn� �����o��<�w  v(�ǎ���麈�⑏VY��Jm�r0�zfT��     ��ɨ��V/l�ӳy��C``��`m��ε��v ��/����J�����x�}]���,��ͭX��k�eZs    �iT�u��V[�ʾ� �A����[������w  �A�8�2#�
��������+��>p�T�d�ˣq�)�    ��*�j��f��L�R�i�ˣ��A���u��r�o�� �o��kJ���OT�s�[>p��|�msX'�"�-     5�����yr�H��p(�r;ʝ�l������}�  ��)�ē%w�(�bs+�����
�\����(W����"��    WY��Ug6����m�Cc�½,���bq����v �H��I���t;�����3�*���Lg9Nb=3ʚ;    �1�Q��V�_�3۳���A���r��y��moz�u�}�  �[���F�    IDAT���Qr�?�EĻ��#�,e���"ss+���Xji�    �����ōv��j;����N�pr����;��� P
� ��A�hJ���*�#���ኮSr���Ory4�ښ�^    �#'����/l���$���\��������n�������s  ����Bk�����~����M��yv�̭a���e�    �Ɍ����6�U]�"�I�N���Nt������;  OO��i��侟�_���]<qQɝg���5�I���Κ;    �aV�U-]܈���`��4��ɬ�z�����z; �����Zs�F���>��gUr�ٛϳm��b^��i�    ��Ɍ�l׉����"Ͷá�3"掕������U�S��;  �L����ƺ�C���XD���.>��L:�NU�h�+�i��%w    �C���ڥ�:;V�N\��;#bpP�v���v��9�;  �L��2��#���GU��>Y���*�·γ�=���(׫"}a    � ˨�v�����g�f��A+�v�k�.�����~��  |{
� �I�}��٣����h�C�����(W��X��    p�TDVnnՙ�Q[��m��h�*2]�q�e��o�~s�1  �<
� W`��^���_���]<qч�s�=��p����    ����k�yf{��]�!���ap����ퟟ���s  py \�̈�A�~��M"���.>�:�͢���ڶ5w    �^Uums+�ll֬��aU��
��4�پs  p������a�~�/"x_�|�L��Mg9�b�;    �~ʬZ�k��F;m�3�v����}�}����  \> ρC����OU�����\)��f�e��6�ղ5w    ��W���(N_�j'����a�_/������A�M7����s  pe���A�hiT|?}����;����C�ʘL��p�Qe�    `/|m��b;3��A�q�g/��|�u�I���r���o�����;  WF�`�V�%��ks+������_RH�[,2�F�6�k�     ���k�[q��V;Q��Y��r;+KUל��s  p��1vIs������������s�1�Υ�(֣*=S     �AV����������Lv�B9�n�e�����>�w  ����]d�`�UE|����b6WH�[t�[��:�Ɗ5w    �+UUms+�ll��j;z;o�v�Ჾ�-�|���;  ώ�;�.Sr�ǣ�U�s_�[J���Y��\�.��    \����b��KV������I8|�e�;o��<�w  ��
 {`���E���K�����c_���;]�p���    �QED���:�1l�}�vǠU�r;�Й���ݩ���  <{
� {$3biPa�yM�#���.>��*����Y�F��-��LEw    �'eFM�k���yz6o�w`7�r;���N�ǻ��y�9  x����`��g�UE|���|o�l�������$WƓZk�]��    ��������:�5�F��Q���r�;�}�7~��7�� ��F�`ZEs��>����{g�6���=�y��a�X�k�2��    �OVM����ک��j;�mP�~�9�2"�i��}�  �Sp�'����6�"~�.>�E%wvOU�h�+�q�eFez�    �c ����.m���d��w`��uZy��-7���/�t���� ��N�`e~����������UU���=�E��a���d�    8ں��S6���¾3%��u�a�4������w  v��;�>�)����x���T����鶒;��*c<��Ѹ֭�    GNV-�Z�p���LK}�vנ��aw�ͳ��nx��  �K��ܻ�����x�[����>|v�|�rs+�g۱l�    8�**�����DWF����Tn�X[��uKß�;  �G��'�K�
c��o4������اʇ�.˘l��p��U�-S�    8|rQ�Y�����L�m�w`we�q)�sT|�m����w��s  �{�z6XF�CU�?Z�Tu�o��]�p���I���.��    �AFU���F;�5�FXm��&�����;	쎳�������?�w  v�R� �y�_�Ex�����g+�P�ju���zv�l�m>�k�1[^�YW�\    T�q�M�}'�FfŠ����Ȉ���_�;  �O�
��h́R_.mD��}]|����}U�I.ǱU��9    ���-�Z�p)�*��QUє�9�n�~��7�¹�w  v��;�b5�?�Y�����UU) ���̭Q�mOk�et}�    �����K[�ً�\�Q����%˃�����}�  `o8� 8`vJ�]y�ǟ~���+�# 셌���\�h-S�    �Y5����yf{6pgG�θVK�^=��<�௾醇�� ��pXp eF鰩O\�x˽]|�KJ��E9��h\kYQ�-    �~Ȩ���Kyvc��"��D����p�ȑt�j7���;  {G�� �Ƣ�����=����.�hU�? ��|�mk�y,�k�    ����ԅ�vr�H�v8����v�v��;���w?��s�� ��Qp8�Z�h-B�}�UE|�So{�b2��ިȘLry8���k�    �����X>)�N&m��8��ʬ'��w�מ�o��/��}�  `o)�-w^!H?��x�ﾣ�Ǿ�x��Yt�[�\�Nk�EtiV    x.2����f����WUi��Q�s��z��+3�ۦ���  �=uI�C"�~ �P��i������I��m����6Gqb>������    8�*&�����yz6o���۹Gl��q��<�ԯ�ӫ�m�9  �{3 ����;��*��\�滛L���;U�I.Ǳ�2�   �o�et�y����g���r��v8��r<��tݍ׍�J�9  �
� �Lf�,08���c_���wt�ů(����̭a��&��2�t:    <�������8���֫��8ȬX��p,����߾��n���s  �?�������a2���=]<�Ѫ*��<��N�f�r˰�    <�"�j<�N���N�������1�AsE��p��|������w  ���Cl��*BɽU��T���_1�C`oUeL�mi8���*[��;    g�l^��/��d��w`�Z<9�G_fƝ�L~��  �/w�C.�����/�_���{����!��]�p�VG�Zk]��    ��̨�llֹ���zE�	�G�V��j���'���vͿ�;  �K��ȌX8���l����x�Vu��1{o>϶�'f�Xn��   �ȫȨ�ǩ�کټi��1�Q1h��@��Օ�n�v�'�� ��[�;  �g�*�.�+g�}���*��X���VgN��a�eL��4��`u�fKK1��   ����f�8���k����o����;�?�����O�� ��� pĴ��\���昺��{�u��[rg,���$WF�Xˊ���   �Q�2��\��s[M������1u������3��  �C���ƊCŏ��/}���6�G<�H�z�l�l���/�m�b}��-�K�)   ��)�*+7Fu���vj�H�pZESn���x���w  ���w  �Ff�`�2�eߙy�t�C�b��;���g�V<~��/ou�զu���X��c��R����w�K�    phd�dZWGm�b;W��s��ѝ7M��������  �G�	�ˈ�V�Yq�-�?�-N��;��5�x�]|��UU����.r4ɕ�8֫"[f�w&    �dt�E-_��熣�r;S;ojVn�Z_],n�����s  �/w�c sg��ܙȿ�c-n|�C��V�OV�������;�g���ru4��̨L�    $-��n��F���ٮ��>O-+���� �؋o����u'�;  �Rp8&2#ZV�,W���d���N�����o����<�d���/�mn����VZF��_    �_Y�1�36'�����A�h��=��������/���}�  �
� �IF��Y����|��[,�u��f���w��j6Wtg?eLgm�9��y-����D    p�TDVM���'.��9��c�b�*��p�-��u���� ����w  ���k+n�%���V�=����T�ϟ=Z����W���uW�e�MU�x�ۭ��Vc{0�EW��    {�et�Y���jk��̝r;q�͓���ξ��  NM ��̝��=���nq����}�E���.>�ɪk��E�9��h�-Ӣ;    쁖�u]-]؈s[���y�^Sn��;}r���[�?�w  w�c,s��le��59�/�'���OU�x��������E�ְ�M���2�L�!    슬����՝���N�N၈A�h���/�m�˯�M���  pp(�w�2"��eߙ�ʗ�XZ�;����W+~�]|����c{���a���by�螞E    x62*[�x\'�_lg�g��@D쬶;~�ox���O��MW�f�9  8X� �;k�����W�8s��P��l������홢;��*c2ͥ�Q�/�5hY]ߙ    �𨈬n:�N<~>΍&��Cf��@�������/ZzE�9  8x���̈��NF��[�z�7���s_����w�ǔ��G�E�&�2�zUD�Tt   �g�2�ټV/\̫�F��g����v�ہ?'[�u����ם|��(  <
� |�'K�˃�W�p�˾;#���b<����]���Ew��XdG�6�ZfT�g    �IF�u�ta��mlֻr�|àU4���-n�n�����s���  LK} � ʝ5��ʗޕq�d�{����Y����O��+OT�����j�?�c�ȶ��+˵X]�툈*�#    �XVUK[�8�=k�ŀo�Q�Z�����Tu�uÿ�w  .- <�̈̊[o���iq�9'p}�F���.>��*��g{��ͭXߞ�J��2��    p�dTD��Q�>��Rn�C���r;<�>zϯ�醇�� ����g��2��z�_�ь���$�/U�d���_����N�2��6�Ɖ٬��   82*3j<�N>q���N۠�H���ZŠ92��s����_�}�}�  �`Sp��ˈ�"���;�/o���w����o���?�LU��;��ʘLsik��y-}g   ��WY5�vW=~!΍&���N��ك���4�z�]ӟ�;  ��; �-s畊w���W�8{��D��|��o����W�E�&��5��"Z����    �]E�n�=�����h4X��S�[e�۽���o�<��?s��� �����ɌhYq�d�O����:���W���ݷw��o͝�-�,�Ǳ^]��;    �U�X,�|�b�zs��W9�Z�z���$p��=Ӎϵ�?�w  w �ܓ%��A�+~0�?�bi�w��k��x��+����Dɝ�-��q��Ʊ^�2�   8v�����Kq��ͼjѩ�Og��ޚ��v���ܾ�����y�Y  8�xv2"��+�5�'~�ũ��u�}��;k����;�|�9��dZ�-��    ����ڥKu�����|��<���j�co�/�y������w  w ��̝C�sg"_�����̿O۳��>�Ž�[s�؞�`c+NL��Ҳ�   882��.�Fu���vz�h�O�gԾ^n�;	g�ZL_�c'��  .h x�2w��?�C/��W ��+~ǚ;J���6�yb{;�-�   Ч����ѸN��883��Aߙ��n��ޚ�m�\�q��^����� ��E��ݑ�""*_|g�_yE�k}�:޾�����VM���U��\�Ɖ�,�[D���
   �~y��>��'.���I[�;p���W�gÕ����������}�  ��Qp`W}m���k*_��7]���}{����}G����;GU�d���{�<h�Pt   `�dTf�xܝ|�b�Oہ�Ӿ^n�;	.'���U��;  ���; �/#ZF��T���d��ӡ_�&ӈ��⾇��Ew���ɴ-ml�U��    캌�5���/���d����<�Vњ#k�R/y��~�u�.�� ��i��  Q���^U�һ"�;��]��b<�;����/U|����Vw�����k����ZZ]���RnWfV��   �+�Q��q]5��/�JdV��������Ϳp�_�� ���I {*�,�_m��xM���wط�Y�C����V���s������(N��4Ȱ�   ��˨̪����qn4n+ہ+ѲbД���:u�b�Ew�+�� �����ˌh��R��?�����h�Ի/<V�;o����*Sѝ��*c<���Q��[*�   ��2*��ɴ;�ą<7ہ+6h�9��g+#�wN~��^w�b�Y  8����-"���wF�ď�8uUߡ��"��኷>P�9Tr�����$���qb>�,�   ��2�=Yl?1�����\�̊A���3<7/x��C��ƫ��s  p�)������~���׾���h8��x�[����>U������"Ǔ��5��y�   ���j-�����_+���f�ʵV1h�xNΜ��s��}�  �hPp`�eDˊ�A�+_���l���w(拈~������Rr�`Zt��I�l��D����   p���b���fs8XSl���b{s���� ��wN��׿��Q�Y  8��GFd�y���V���-�>�w(""��D�[������2��\�ŉ��[�Tt   8�2�eu���nȬXT8V��qǭ�����?��� ��C��^eF��8u�򯽺�K�J��< O�����.��������2Ǔ��5��y-��N�   �ɨ��f�����j�v�jmg��gO��׶ӯ�;  G��; �{��>h�?�ݙ����+}�""�¥�{����U���\�.r<���(�g�ni�a�   �0˨̪ɴ��y��b;�eTZ��1��A�K_����;�}g �hY�;  DDDF�\MT�rC�k_����W|�q��}�����T<�������n�1�"q`-��Ť-O��WWk����]E+��  �K��5 {+3*"j<��F��R_���Ί5S�+ײ�Ym�]w��?��9��}�  ��Qp�@��Y�8��W^���OE|��+���d�&�=�ŭ7f���g��)�spUeL&�<����J�W�s�"��s  �Vf7���}� �hʬ����ck�O�S��\�A���O�}ϻfv�_�ʙ��w  �&w ��hQU�һ2n�6�]��bs�w0"">���e������� Ca���*c2ͥ鴖VVb��R���   pPdET��p9F�PAvKf��j;�����}���s  pt�� ����ye�5�*������}ԃb{��W���*6��8�*2�۹���'����"�'_w   �>ˌx��-�9����_~b=����.j��w�ŋ���_�'g?�w  �.� l��m����W�<����`�E����x������yq�K�##�*6]�t���N�,�bm5�]�/~   샳�#�����RL�[Tt�O+��#�����{���'���_:�_�� ��M���/���t��f�;����wq�RϹ����"�C\��W��hu�9%w���Y�gube��,�Gt�G    {�k"�})ΝY����l�Z�~o�k��x�C]��}����j;쩓k������  }
� �gOE��W���?���OT�����F����ŝ�f����X]Qt�0��E�X���vVT��    �Ufčϋx�m+q��R���o��֌kζ��}]\�����aW1hV�a�eD|�G���o��}g ��Sp�pɈ�U���⌛��z�.6��FDDUħ?W��c���Y/yAF��;��׊4�Z]��A�]�N   p�d�x�M-^���X[]�E����?�������-�`ş=���@�    IDAT
\�̊��&���?��������s  p<X��P��y���*_�c-��'��t;���x��6�m��|�9���(NT9h�H�?    ��� �;2^���;_���˱�.��vy)�/�x��f4���3�)��r;쇳�����S/�;  Ǉw ������R�}�M�g=��.��}�k��x�[�x��^����5w��"s8��A���n����]D�V   �o�����Z<���DUF���2^�����T<��.Ɠ�L
������A�K_<����]'�� �o�8�2�l�V<����m��?�x�1��E�E|�S�~�������땃9\]�bҖ�Y˫+5_Y��HEw   �;�q�������jU��>��]��j���+����^`Gˊ��� ��;�o��9��}�  �x�r? ��̝C͵����?�-�|��@�F���.�{�j4ޭk.�?U�i[�؊�i����ev}�   �o��D��w/ū~x-n�n-ݓ��]vb=㯾2�/�3 T�r;췛�7{�_�ʹ���  ?� �St���붌�i��G*���� ���*�����zQ���(#�
6�M��,۳8��T���-2+���Š�NI`�U�Um�w  8�2#n|^��.����1_d��ῲ33^�]�NW<��.���gIEf�@���ɵ�?����;  Ǔ�; GNfDFũ��?����}*��\�Bzp��x��P����uW+�s8�晳�`ii����"ڠ�*#.���-�-�ڢ�<"��  ��� ��g�q�r,-/Ţ۟b��[3Νiq��]ll��?�CŠEd*��~ˈx�F�t�?��s}g �xRp�hʈ���K�ʸ�ڬq�qМ������֬��=�+��N�E���ŠU��,b0记�   p���F���ݼ�躌E�#"gOg��[������+e�e�z���O>��7]��}�  ��Rp�H�ښ�5�"��kZ}��+>��U�3��*�ӟ���+��;���E���w��u����{�A�F �IQ�&;v���q�N���=K�T������LZ.;v:�[���L�K��z���{*����^'��rǶ,[�J\�E�A���X�r�g�8�D9�D� �]��*e[���!�{��92�
F}J�iq��\���
Bw     P_�:�];m(���X[�ł��?&�8+=�o�Q���@�z:�}����=   ��; ��ls7s{�id��w��Z\�{0ܭZ��?�:���w�F��ѴT*�ʮ���X\}o7_�     ���I��]c�z�
�VUҷ����.�?a��4⩨%�z��`�
�9ErT,D�5Q����j޳   ����  `��I�\��>�A;�8"�E��ҟ�e�7�t_\+ZP��M�J��bQ�r"w6    ��Q,H��G?Т�<�Y�m�T�&us(��+�ģA�����.�g���hf.�X�?��X�_�=
   ��= ���������(~$�9p��	*8|�e�������-�k7y�m-��#�>�J
R_�Ɍ�cԷM�j�4��aM�R4�+ҝE��˓c �C�IE
5� ꃙ�`馼�  <���ҡ�A�8Ԣ���%�^��ołl�Xv�r�v�� x�l%l��r76R:�{_�����    $���   l������=f62�ɣ�K�ԥ��R��~���Y���|� �;�_���҂Bٵ�5�}�J�D�D�9�\�Z     ֞�4�k�5���;Q�ZP�A>j&{��@��w�FU�yO�^s��y(P:�b����=y�   �"p 4/�O7��>�~�ū�O�*��?l����5>b��æͭ���M�r�r9Q��wg�=�A���^H53ǃ     ���Ei|�41RT�%Q�T��=���uu�ɨ�;yO�G1s˾��b�~p����ا�f�   XE� hzf�6��!��^��ײ�]�']����g
F���*ՠJ5��D�E��a�5#�����dT�yO	     �M�VibG��PA�J����ͻ�e��h��<�p�s^��da;[ہbAv-�����qޣ    wK� @}��}�C�n?���w�D�o�$�T(��G̺;M�S��A^��H�K�oHg/�6o2uw�����T�UӠ-�M�C��H�Bb��#�I p�ܓ����2�,ݔ� ��L��gz��D���h��1�{s�� ۹ôi�49%9--�;�+	��@�ݾt�������   �alp `�J��6����(���N�7�;L]��h1��K�J�b�upO�}A���]L53�u	     ���ŴsD)����J%�T�{�|���O��;̿�T�r)f��v�VulM��t�3�9   �7B� �3)ȵy��#�7]�j������jյ��g����yش������T��ʕ�b!j|$�Ĩ�֌�ʥ��WS��    �ĺ;�]���oK��DiT��=Um��'��G�?���4�-�����f��jM11߻k�S���-��   x#�  ��^�k�6�z�.���|�u���	�D��R�U�A!��ۢ�}�tho���Q�.F-.q}    �$A�n�3��mKA�JP��Q؛��*���̏�^<�
��9[ہ�w�ҿ��gz����    ~w  ���6�V��׃RY��s�Sg]�	>4@���i���TNT,��7a�74uS:s!յQ�s#     N�V����ႤD�j�2�o��렩����G��ռ���+[ہZ6��t�_��d�s    o�� ��b�*p�ktHls���ҟ};j�v��1m�B���.�+�ʕDI�����/�/$:)��Q�2�)     ꙙ4؟mk����*U�������+�_|/jv.�i����v���oMˣ[ߕ�   �[!p �^�$mnu��׉K���S��{��3Bw4�45-�������>��W]�.����     �d��l[��p�$)�\Z.�=U�ho����iץ��� ���@}(&�Ɩ���??8��,   �[!p ��x�6wc�{HS��Iי�w
�gL��ј�M�J�R%Q!���5M�v�r)��dT��=%     x#���w���$*WUӠj�{��T,�}�����g_t9G��}ak;P',����?���{�(�Q   �{��= ���������(~$�9p��	*�y��J�^(��G̺;M�SN8ZêU����eW{����_hl�M�jP5��j�1$�K�e�iyYl}�Tܓ��� < 3��My� �fs�i�X�#�c��B��J5�;�W�z͆LW���ռ��ɕWyO�^�-���/u}8�9   �{�w  ��ls�9ׅ+l*�e��ҟ'j���#GL]��hl1�J�D�r�B!j�H�]�A�f�mu���J�	    ��2��{L�Ƃ�W��W�J�'kN���O<���\7�9��J\f�Z�EWg\z���#y�   �lp������}ܵ�}lج��t���¶��vgAz�םi[������/FS��(M��l�vl�v�%ں%hi����a�� �����nk�F�*�*W���TފٞqS���ͼ�j��+I\�%�-����W����d޳    o� Xwms�&�ُ�����Ĥf�Kg/�.\u�k~x�)�;_MK����R��j玨�Ѡ[3�Vw     �X��@��XPoWPee[;4�I�����������x[ہ�c�L,��/|��O�   x�� XK&�Z�n�6�gBf��o�Z��?�:{������G$wBw4>w�\IT�$JWG[�w��Ot�J��˩f�xh    ��h�j�946�D�J��2GN�`|D����'����=��l[{8#���h��o�j�/�=   p?� Xf�6����|4�Kg\Ͻ�1���f�,J�z*��i�#G������<�Դ�de��DM��v��n�H�/G]�LU��=%     ���H#ۃv���̢�J5��^w��e����~�u�*q/��+	bk;P�������w�=   p�� X/������#���g\7nq\�n�r��o������������]�T���Ip��E��!�ȁ�+�]�/Eݸ�\�     xUw�ibG��� W�J%ha�#�zW,�}������/�������Ա-�����k�v+�  @�"p `�e�ܥ��������MO�ل\&�\�g�=���8hj�D��FSZJT*%J
Q�ۢF�LK�.]�:w1jq�]    ��Ժɴcȴs$h�l[�r9�=֘�l������[OE--�=����ԻB0߷g�_����y�   <w  6�J�.w�3�ms�޳���ڶ�K/��:wɵ����L�����%U�A�jP�b!j߄�o"h��KQW�"[�     �L��	�5mJc��}q��F7�+�ģ��x�uc�s]4�`���v��Y��]����~ޣ    �� ��dR������?&]��ɣQ�Ky��R�J/�t�=�:r�|�I"tG��T*'*�������~�R)��+��WR���     �Xڷ��GLcÉ�Šr%hq�m��fs��o|����K��q���`r��alp��?�B���   �Z p `��ls7I���~�c��9�:}��׼�e�{G]'N���P�ۉ�Ѽ�iP5
�*\{v��;a�=+]�uq2�\��    �OŢ424>��T�U��*�yO�<�����@����DUӼ'�_�@�4����Ү���    �
�;  y1)��Rt��w�v���h��|ރ�^��K�|2����=�z	�Ѽ���S�TH�:ڢ�yHz�@�Դ�����SQ1�=)     o�L��	1m�U*AK���v���������f��x{�\I lŦ�ǽ��?����   �� ���e� �}�����:v�	A���ۮ��-׎!��<djo#tGs[��n&����T����r�KW]���=��3    @m��0���
�lS{��,�L{��?��O�.]�����,p�̤�{J_��g{��{   `-� P,;�*�ۑ���P�'��n�␹^\��<�6�C��[���ܵ����\�B�=�A��˓Q�D-.q�    䣥(&6uwU�A�j�r5��PO�٣�7?qV���.�5*�+��h8��K����;���   �Z#p ���$uw���G��]4�����Rރ�^�K�/�.M���2x���H��h*��ʉ��ڲ9��^���k7��WS]���yO
    htI��o6m�Jc�r%ha�#�?w��	SW���>繨-�,l7.s@��V��;���Ѽ�    ��;  �Ɣ��s�4�=�s'\'ϰ��^��t�e���\�w��k*�IJ�)-%*�%I�@o���Z-hr*��ըk7"�;    ����4��
*$a%jy��3�/��G�?���4�ț+	�_�@#�j�.?�����    ��;  �ʤ`RK��æ]��OuM��0�^T�ҋ']�Ϲ�3?�����$�TM��i���XpJ;�L��DW��.\����    P��l6���G��l�TU�A�Jޓ��mn�}�C�G�gg���s�B��hT�-1N��~��?��V޳    �� �g��B��K�7?b~���K�
��F�,=�m�?r0��1I"tV���S��W��sG��h����dԥ�Qwy(    xsł�}[�ذi�'��fQ��G1�P������'�FU�y��fa���lmW0ׁ]K��7~��/�   XO�  �[����OH����9�:{�C�z��$=�L��w
>6,��wK�)-'*����[��+ړ�֬���,v/���    2fROW���it(ȕmk�CԎ����v����f����B�h`�����/�|5�Q   ��F� @���}s��_{�i�������H������^To������o��UӠe������T=]A��]�r]�����JӼ'    䡣�4646T,U�AK� �NԒ�6�O8���4�W'֚�L
�M*@3\8�ۏw}2�9   ��@� @�Y��M��>��|4��W\G_t^u[g�o���/]����<h����Fܥr%�\	
�*\�R�*��&��.MFM݌Jc��    �Ӧӎ!�������J%���*���v�G?`��)鹗\N�5�J�dlm�Bog���Ň�   �(�  �+�6�'�´c��{Ϲ�\�0��\����r����!� �;�#E7�+����UL�F�K�ær���SQW�E]���   �!��������D1Ͷ�/,q����.;�״���[OE--�=�Y0���h[Z=}x�����Z�{   `�� P�,;�n�*��LW��?�l�����Դ�?~˵}��݇M=�<� �L��RLT�$J��P���G^�_�ٌ    u&	�@�i�����\A�J���Q�ze�x4�O�nLs`���e+��K!�4���C�ʿ��O��{   `#� � �$�kdP��'�{�u줳��MN���g��{��	݁��FSZNT*�p����r�uy2���;    �*3���4>48$%�V������ln�}�C�G�K/���Ɍ���������?����   �h�  4������~����=뚜�лMN���_�Ɔ��y���F�܋�c�B�R��3�g��;�+�\����=˵    ���m3YȢ�R9�=���]M���O���y����
&��9Ќv�.?�[�����   ��;  hu�{G��'��������E--�=�.w��eׅ+���G�ڶ����U� +II���oWԾ]E�Y��LF]��jf���    $��'hdд}���$�T�J�v4��;dݝ������;yO�Zb�
�9��P_������    �B� @�Z��.w��!����S��m@u�]:{�u�k�����-�y��+�]��I�$j�T�w��MugI�r-���fwbw    X[�D�4�Y�T��ՠJ5��|uu�>�h�o��ui�C�fg�mm7�khV]qil���=   �'w  �e݋�vd��k4��]�/s8^�ܥ��]g/�v�����R�T���G�0��Y�����dԭ�H�    ����4�o0m��e�b�r�Z���G?`~�����}sr� �v���n���ѥ�|��=��   ��;  �¤`R�V��״w��������{0܏���\v�5x�i+�;�>vwW릨=�Q��Z\\��~��    �Ŗͦ�m�����.S��k�D��w��	SW���~�r)1\fY�n��M����Z�̗��;y�   �� �&c&�\�d��h�S���{�U��=�G��F�3\��G���_�J�^��}Ӧ���=;-�
����r-�ƭ��    jCW�i�@��6SW�)�YԾ�D�܏�~�'>��']7o󫨑���vck;��L��݋���?���y�   �w  ��eeIp�?!M���I��3���^�Kg/��]t���󠩽���_���.))D�Q���т�Uij�u�Z���Q�j�   ��1ˢ�����!S�֠4�>0<��h[Ze���ϼ(�8͡m#
����3Z>�[�����   ��  43��I�Z�9l�=j��s��i�땻t�������G���%U�A���=�*��\C�U�]�u�z��T�    R�H�AC�LCۂZ�R�f�C���JE
!�ƛ��+X��������J�{�   �%�  @f�+P{�d����+������d�_�ҹ��W.�F��y���A�<(�TM��io��B!jx�4<�(Ƃ�g\W�E]�����J    ����E��LÃAI�rOD���RY����Ӯj��4X+&W�Y< ���.�_ޝ�   @�!p  �2��ncC��`�c/�^<�Jy�R�ܥK����\c��G�:�	݁���/��$qQ�=��{��Ht{�u��    IDAT�zԵQ3s<�   P��l6dQ�@�I2UW6�/�8R ��¢��)י�����J�����X=����}�>�Y   �ZC�  ^ϲ�=1�#�M�F͏��:���z�.���p%����~So7�;���Ԕ���KI�'QݝQ�]A��&ZX��nFMNE]�yP   �ft����gQ{_�)z�/.������,�_<�:}���6�\����TT<|`���c}��   �E�  ��eeڷ�>�^i�D𧞋���{2<�Ս�&]�������km5vW9Q�B��5jbԴsGAժt�kr*����R��    6N�H�]A۷�l3m�,Řmi_X�w �of^��)׹K���,ۍ�)�7�uhO�7���   �U�  �M�I&i���g~"��s��^r�+yO�55������J����Z��T��ʕDfR!�*������%z�D�3�k+���O�   ��M-�m�٦��~S� �+Q���@\l�۳�c���-�k���\!d�; �!ڿs�����;���(   @-#p  om%r7��%�	��K�2�Q���=]��������]�T���$%IT������	zh_��y�䍨k7\ӷ#�Y    ���ô} h�@PO�䒪iP��\y�4��i��'\�S��7WB���ޱ��o?��ɼ�    j�;  �w+���Mn?�N�О��w��̡}#�5#=����}�w�$Bw`������(	�B!��-��#h߄�\��ߌ�6u�\�z   �GKi�7h�?h��i���R�4hq9(���y�:%�kj���F���xk�*7��W:ޑ�   @= p  o�I���v��״o��/Dݚ�{0���9�/��q��>��c�`���zK�)-'*)Q�BU(D��F�
�Q�=뚜��v#jv��h    �ڶ������7���4��-,��sK��L~�t�k�67��������Q]<r��/�9   �zA�  dr��>����HO�ug1�ɰ���u�p�up��ޝ�BB�l�M嘨\Id�Wc��nWowС�����k7��߈����T�   �FH���V�vSG�IA�jPZ
|�Qt����^v���{�3W0�qR
�m�+����ا��*
   �G�  �������Ɔ�����Ϻ��tU*y����,=����}���6mj!t6��T�U�A&)$�v��MQ���;���7o��ߌ�v3jn��   h$�[�ՠ}�/�Xp���ՠ��4�6�[�*?����i��r��`=�\!d�; ܫME�vW��/v�Ky�   �w  �6,��^0���H{ǃ?�u�5�A�+ұ���]�F��gj�B�l$����4MTR�`�$q
�m����':�mw���mw/�#   ����ni7m���0I�4��AwM�ܒ�`�$���s,�h\����}(&��>���t���g   ��;  X[&�6��=rXڿ3���]�/s��(�Tz����A���z�	݁<D7Ū�R��DIUH\���mww�f�\S�QS7]7nE>x   Ԡ�M���,h���Rty4UR����΢���,lOӼ��z	�������?��g�~;�Y   �zD�  օ�lt�hw��{��;�?�Bԭټ'�Zq�.M�.M�z��7�J���@^�4(M�R����ITO���+h߄�T�nLGMM��݈ZZ�!-   ��$�z���L�A=]li���Y��Ӯs�xse�r�eq;Wa �ł��Z�O_������(   @�"p  ��,�R�}��?������,�=��Դ�Ͽ����>6,I<����v� ��j��R�2�l7�'��wM��6�߼�:   ���vӶ��m���S�H�j�-�@-3�_�.�x�u�U{#3�B���� ���~�]?��   @=#p  �o%r���K#����u;�T�k�֌����ڷJ���3�@�Ԃ45�i�����^���puw��N�Fi�V�OMG�̱�   x--��^�`_ж~����-�j�h�Ėv���+��OE��͔���Z(_�'_mG�s    ���  l��н��=�G�;�����g(����Գ��^r��m���u�Zq�vw�W1�J��m��@_���\�nLGMM��nF�Y�b   ��$H��A}��ޠ����v1��)[ځzQM�ϻN�v�D��\	a;�5��U�?�maw�s    ������U�@0)������ai�x�g^p]��C�FS*K/w�xҵs�th�����@-q���]Jd&%!�Pp��F��������]ӷ��}r*j��u   ��L���b��ޠ�)I$��jZ.���`?P'�K�S�d9J弧�z�
�4���і��-?���up!�Y   �F@]�m��7.m~�r��77u�=����D�[�ޣ��K���G_t]��C�Ɠ�o�L�f:�۴}�KP����UH�
�()�f�K��i��[Q7oEU�($jT��	y
 < ��$�ܑ�@�ڶ���z����%;�H��Z�6�G��'�3�^v]�&�a;�����G����_�z&�Y   �F�	+����o\�9}���͙dk޳���nx�E��t��/Dݞ�{(����d��Sڷ+hbTJ�)�^��*��I%�����9��k�V����� �6�Ѭ6���{V��>S��ܕƠjTMM1r_�3��k��Ӯ�)b�f�e�2.� �Ц��:t�{���?�{   ��p��|�_L�~�ٶ�擖�g��#pG�Y	�%�W�g�E��2��W�m�,�eڳ��R�r����Z�\���(ݚuݘ��1�5�Ƽ'F�"p��A��fQ,J}�A�A������d1ګA{����p��T~���i������F0�=�I 4�bb~����~�z���,   @��6�}���̾���o/.%I޳�G#pG�Z	�c4?sQz�弇��{�w����1Ӂ]���\��zd&%!�PpBT��dJSizf%x��=	ޱA�`m��QR_OP_OP���C
!{�\5�VMir<umiY~���9W����`r��� �ւ��[��o�J�g�   hD�C �����z�xǿ*U��E5��u�%w����8�:v�U��=޾��W�Icæ��L�\��z̕�lw/$QfY$�ҫ���[Q7o�lxO���� ��;E!�z�����=Aݝ��i�E�ij��~+��ݞ��t�u���A�&A�`�����-��_��ο��,   @��t��կO���':~�\�厵��å�R�b��i׉�NYW�
���MM쐒�KP��ޓ�e�r7I&w�̜kz�5}+jj:����F�`m��^%����ם}���ǔ$�@#3�ONI'θ._s���4\	a;��o���������=   ��8��&~�k��8zb��OyTs��pVB��e�N�N��U}x�� 6�J{w��M�Z7qI�j��������]��sݼ�y;��^.s���!p��A��zQ,d�{�M}=A=]R���=��U�v�QUS����g\sw�)�+� ���������   ht��X3������S[��������a��4wG��qׅ+��mm��$��GLv�z������UH\�ʆ��\ѥlû4�u�kz%x_\�{C� k���jS��o%f��6uuH!HM�hJӠjj+oЈ��'ϸ�\tUxXS!l�����&��ou�=   �8�����㷾}�\�\&�
w4:�l��m�3/�����S�־"���B��;$3.s@#2��U(��WX���L�%���ׂ�۳Q1�<4j�; �wԊ�MY�����e������n���vv�v���'���_a�E3
�2sq,`�l�-ߚ�����gL   ������_~u�������w4�\ك�k7�O��5��Px���
ڶH�&L{v�Z�\�F���{\�����*�Z	ާo�n�DU�yO�Z@� k��yi�j����1���ڶ�L���WSSJ�4�J�u�b��}�N��`����v�� 6R_Wu�=�,�=��n�>   �{ k�ܓ?�ܝK����=��dVG���Kҳǣ�y�U#ֿ2(�����L]\��f`&%IT!�B�J��w�,l2���o�D�3��EV�5#w X��I��:�z�M�]��nS�&��Jc��=MMilk���ש��3]��qh2f���=�I 4����һ��~�Sm��   h& X��ƥ�Ǯv]�:�ғ�,͎�Mi%t����e������5z�ݦ�L�#R\�f����lxO�ו�l�P�J�u{�u�v��\��+yO��F� k���X��;����;�О$هc�6�gA;�v@srMNI�ϻ.\�>�B������@^:ڪ��U�;O�=   �l8
 �n��W��^�8u��-�Y��;��{��=�[Z��1��	Ӗ�\
�fd�Wc�B�mz϶�K�[����}5x��s��6w X�X[��J���mjo�TD�"�t%h���F�����e����ٹ7�;��j؞mn�<l�+�8P���뙼g   �'� ��7�٥᧏��<=[؜�,͊���B�3��G-.�=T�ɷLA6��e���43S��=ޣB��8�lӻ�J�uk�uk6f�ϰ����� p�۵���������%��Hr)����i��/���yשs�3]�7��znTfN� w���>���<��gy�   4+� ��������>?s'l�{�fD�܅�=G��z��K�7�sD*jf, 9
��I�W����K��r����l|u�;�{� p��A��7c&����:Lݝ�v�����w_	�cP55�Ƚ�׸��\�N�q]�q�oԢ~n4�� jŦ��#{��/����   hf�"�_�ݫ�~�D�w�,�b޳4w��p��R��r�C5��	�W���Ӂݦ���@�l%x/WX��%�n˻�k~�u{v5|w��F�1���#��� p��Z7��;�
�{��,w�=�W��{�U4��e�ً����ŷ�OSA7
�v ��������g�� �Y   �fG�`�|�����w�n����$�{�fB�����=M�_>�:vҵD�Nj/p_e&o3�0�J��Y���+	�_K.��fJ�kv%v�=u{�5�^�b=��� po^�D����2�t�z�L[6Kr)�)��4JSS���? 5�u��t�����_���w&W�� jG1�?�w�_�垯�=    � �׾q�g�=���.�C�{�fA���6�US����G}[Z��1Ӿ	���u12��F�I��}�|�gאj5��>w�M�y"p��A��B�ڶ�����C��2�b����,l�{Q��.\������[��F��zE��sٿ�;_���O�=   ��� 6ܯ����=}�����5h�o�]���s��N�J�pk�>�Uf�`���n���w&e�WQI�6�K���0���躳���F�sQi����� ��{�1���^�ww���}h/��A{��"x��g\�_q��誮�=ut�1s#lP{�\����ϯ��ο��,    ^C� _�͙�<{r�?�T��7w�>����
����&��i�5f��R�? 91���mx_޳��5z_��>3�my��_� �y��� p�ofRG���3�ٻ:L]R�Hr)�+[��,l������J���%שs�۳���B%]/��2�t`��������g   �z�P��?�G�����-�U#ע�D�< �\R�j~��œ�r%��U��I"����4���@����J�x׫ٳ�=�+���΂4;53����e����� ��{�A�l7u���ww��B��=F#f��nϹ^>�:w�UY�34j�ZG���Y����'~�v=��(    �*N���s�>�/_8���D��w`�Ć���K�]'�n�C�F�X��viטi�8[����6�����ЦwI�T\�+����W7�G�l{���`m�צbA�h�h3u���;��.SY̾�Ǖ�Ng`��uyRz�׵�����ZE��^�]~�����H�s    xc�8 r�����W/���?ļiP������/�r�H��Qc�
�4�#��{� G&e�{��ae�$�M���%Ř��+��gW�-�
$w X+��k�d�l7uu���MݝRۖ�?���=�c��� X{�3�ӯ�^���"��Zc��P �m�p��?���y�   �G��P>��[�♭�-���;�VB�j���׋']��yU�3p�[W��g�41�Vw �+X��nz�W����T����M��;���DB� k��}� �o�6�w�|��0��Jre�j��-� ����+�����l��PQ�_�p6a;���c�|�_�f����    ��8�P3���p��֟�{�FC�����=��g/J/��ZX�{�Z������ѡ,t�&�5�@�����ޓ�E�o���]�w\sw��sQ�4��7 �; ����R��ۂ�;MmRG���Ӕ$���{�f�{��^�����]rU�yO���:of�`�� ���@��h[���[���   ��q��|��3��K��|L�@y��`%t����e��Qsw���4g�ѾU�=f�=n��ڔ? r�m�{m�{����]���|��B���q�/��:�	�`m�?�$���λ��wv�6�HrS���ՠ=��߯`�-�\�.�N�w���=���·�L�� ���@���O��x��qF   �* 5��o���-j�r���W?�c~����ٹ�g��}U7�FM{�MÃlu����Ǖ�=�O�(|_\����;Y_���cx��`m�ߛ$H�m���YĞE���-���A1Ji|�{Bv ��59%�>�x�c������v �l�@������   u��@M��~���_>��=�&�F������5��㮛���z�܁�ݶ�J�V���o�@�0s��W7��+�K��$--���}n���;��Rm��G� k����VC���,b�;d7�b4E�6��i��ݹ5P��\g/d���,�=ͽ���(Yؾ��h �?C}��c?�>B�   ��" Ԭ_���s/���0W�C��h%tw7]�!����t�>{���afҶ>��1�ذ�$��Mf��K!�Wxӏ�+Uם����ʷ�]M7��@� k�Y�$�ڷf{{��V��Bv_��WB�հ jY]�'�3\W�{�I��}��h���7����   �CI��g�Σ�������g_�� ���%1�L�G9n��ݓƉ����c���-2"���GA�"�Ѳ��q*�i�&'I]��/�j۲.�����ݟo�x��A `��.��93�f��������=3���ӹ��[�>w�1�G���v�k�kp�7�JI;�M�w���$N�4��j�ޗޮ>]�-	d�z�V*��j�����YW5\�����h��=�����t�:;T�M���u��am2{H��9MϺ��q;�*�^�J�����u�� �����ć�N׶G�
q�   ��Kƽ  ���d�}�c��gs��9� М̢�Р��ӕI���F/4�,��rY:~&����!��nڷ���ɕD �+tSX5隉�&ɂh�_"�4|eŃ�^S�ii���|AW����%������w @�	)�����.��#����cJ&%�E���졛��єv hV����9���P�q��*��N��5���\���w�   M�-
 odă����'F���^K3b�;И�ݧf��8�:q��Cwj�[e&���0��*%�
4?3W,NO�BxjA�ڏ���>�ݵP���]s���\��N�;�`u4�� �:s��vv��:��.��3PG��i���Tv� h!a�� ;�:w�����Z�� �U��.���'6�ƽ    ��{ M�sO�ѧfN�:���Z��;��������G\'Ϻ�0�U�J��H����Lw�a�0�_%��S���j�����遶$�y��`��8�}!�����+_pU�� �)pORg���5l    IDAT��#�uv��Gq{��^3��C�9���)����0�bK�����@+�4X�����m�=�e!�    X� Mcdă��̱S�;�^K3!p��K.�P4?t�u�X�]�$p_-�=ҝ;L�w�rY�Z��z�ԧ��_��2��w���9�Е/��|P�_����g���y�ܼ{�H� ˵ށ{*�ꝵ���SW��ܒI�a=d_��ޤb ��B1
ڏ�vMNǽ��B�}{���M���{���   �� Medă�٣'�evŽ�fA�4��D�r���i��]����W��4<��;��d��b ��l1�X�����wW���dA�����ժ�|�}!//� ~>/�_�/�y��|v �u��'�{G�ԙS�uWW�)��&�������� �,]�.J�N��]h�g�
���j�� ������@y���OŽ    ���  ��Ȉ
3GO���/�;Фj����Ԩ���PS3q/j%��R2)ݱ%��7o���� i���@��A�)La(��{4��:�+7/]]�_��x m�V� �:��{G.��^��H�)�K�u����]�p�<�Z���n��r�-� 0 �������<P�I�   �� M��}�܁&W�%��қG]c�����z��J���v�a��� n�6��M� pO$,�^�[�0�B�䒹ܮ7^�ª�BѽX���������kS��9�&�fwm�n&e3����n���]9)�5�6}�]o	י� �73�'κf��^M��ؾ1�Y�,W�@ ��6������92��R�k   ���� дFF<�P�9rr4�[L�!w�E�Bwwib�����f�r�q����0��n�e�' �[�J�2W"P����,��P(Wm
�jS�op�d|��
򅂼X���b��4x �$��e2�Μ��í#��3[��̙rY)�5����aMe�G� ��S(�N�s�8Mmǵܯ'��	����������=��   @kb{@S��bi��	"�"pZ�{��-�w=�T�^�;!p���4<dڽôcXJ&�� ��ru
��s&��)�@^�A5����x�$y�����P��� ��������j���� �M"�2Y&-K&LARJ�[2aJ$�DB
Y:)�3R6-�2�lF��ȒI%��ͪ�a�w�0T@� k�Zu�9/�<�:�r�w�\A=6a�@���_�{h{�����Z    ��9 4�Z�~��hn/�����+
ݥb���	סc�b)�U��{�H&�[����� �� ֚�j� Ph�h�� �Ln�"y)��)��������P��KQ _(�K%�B)z�P���b�U,�`	h��,�1eҲLF��ʲiS:�˘e2n��)���R&�e2�����M�
<��u"�,�zF�BMbwc� և���e��Yי�r9�5w[�@;��?���}�Ѯq�   ���*��02��������Lr��;��HE����Ӯ7����^Ե�Q&-��fڵ�4�A�� ����<�
�f^��A"
�Y��n�d�<^��͋EW��8�Pr��H^�r-�/�J%y�$�6�3� ��L�֦�粦lZ��Ȳ�(dO��׳iY&m
nf��p�̯�`�K�ah��e���z��� `�MN�N�q�<�Z(Ľ�fԾU7a;�v6�W��70w����Kq�   �����12������g���;�Fj�{���^;��l��CJ�F�����{�����J�f�̢��6!�M�V{=��VK���G��w
�%�Z5/�\��<��]��E!|-�/�]�y����y��(�@<RIS&#ˤ=��3�D�t:
�;�Q���n� �sV�̰�^��Y��G�z��Y�`����=P�i� �4�\'G��}j&��4����k?K��mm�/�<�=�����Z    �=�| h)##\(N>y�c�{��hO�G�s�7���.y�m�����&��#��fڹ����? 4�ڄG��.݃ �ɢ��f�[ 7�[`����џZΔ��ܼ\v�*楲�R�B�JټX���R�"/U\�j���敊�\az<���I�2S&%�Ԧ�gӺ��2�TZ�IE�z")�jS�Mo���[(s���T��.E���m��n �Ɨ/�N��N�JW&�ޟi%�SyGa��8= ��6o,M����=��ឿ   ��`+@���Je�{G�t��Z�;��ܣ������'\�X�1�f�q��s[4�=�� ڃ+��\���xyԃ]s�b$_�_:�8)�V��^w_����y�ɗ+�J5�_�F�|���T������r��劜�K%��t�-���k�z:�꩔,�6�ӮL��.ˤ��_߮�gBp��ea=Xw7�)t�MW�\�� �Pt�>�:}N�x��}m�z��
)h��M X���*w�T�#�Z)�    X?\Yв~�3�u�T�����	�H�j�{�b~���#��u�sB���̤�M���vl��)�I �M�,��-��&�-����R�~�N��^�_���WkS��Uy���ˮJżXrU*�RE^,F�+�\�ڄ�r��L6�t�+�����T�-�6O'�R)S*eʤ�t�-���YjƂ`q��$ES��o��W���Z��6��
 ��R�u�tj��I��b���A4�  m�T<���{�ȈU�^   ���U -���N���;Qw	� �"
u��gǤ7��.���}$�{+	ixȴs�i�bw �Z�����vɢ_�P^����KR� �d�������zK0}�[�W<�*�B�U*E|��*�啊y�����R�"��\����rżRi�ǡ�jix�w�I��I)�4��R2�LH���J�IW20�SR2)K%���dBA2)K��	����Z��z�MH���R�x�E�U&� �H��:;&�u���
�w�3X-�U���#l���.����zwǽ    ��������&��7�v|$�uą��u�r#wib���Q׉�k9]���U��eȴs�i�0�; �����h���߸�Em�|4i~ɛ���%��j��kW{_(y�,�J�rE
C��*���R9z{�b��^��˥R9:%+���t�l��]����S�boש�� �0���,��	��fq�mfJ��@R2����fQ����dB2�%��L%dfRx$OnA K���%�DP�~.In����hNi4=}��~  X���Mj?w�U�ƽ�v�%x`.8�k��R8��{�{    ��~	����s����ο��$ww ��=���O�sK��_�~�$Q�~Gm�{*�?;    ����.\�N�q�����f�]A�� �kX�;�-|�W��'�    ��	�������ᎏV۬�$p�l����������á�gV�s?�f��    ͬ��.I�c�3�]�b�+�[5_n���:O� �$�������s��{)    �Ge��<u`�7�8���*a�����e��]2�$<����]{#pogɄ�u�i�6��MR��    Ѐ�U�����h/�I퍬y*q3W`�� p3&��=�?��/��͸�   �1P� h;O�������J��r'p���mv���	���J��>�C��8�}۰i�����    �O���,�u�#jo�^�GQ{4�2����ޕ���<���q�   @�&Ж�yi|仇;�-W���	���Z�^��?�z�k~�>�Cx3i�i�6i�6#v    ��R�5vIs�>�T�^n]#�.�Lk��
�w_�߾�L�ߏ{-    	����/\��뇺>Wj�ȝ���r�%�����ҡ㮋W�s���7�4v߱�ԑ�K    �zJe��t����%W�������
r�hb;a; ,_"a~���|�ف��{-    �����/O���_�}�X� w k�]r7����t=y��g�5}=�[M���z���    ܺb�u�B����
øW���%�b���ct `�%������O��b�k   И�n��>�������)�D�kY� ֜G�{�j~rT:t,����>��!ܶ��(v߱���͗    ����]gƢi����2h���w�+�� �+�pp��K/|j��q�   @� I�}��G�����+$�q�e��X7.����'���Μ�OG#p�����m6m�(#�    ��MϺN��F/HSD��a��r�ŉ� �ۓJ��W��O�>�Z    46j ����ϼ���ߜ�K��^�j"pwI.���θm~!�U��d�Ҷͦmæ���d��    �w��	������shG�U�GQ{��JeR>���������^   ��G K|��S{��z�{�Ɏ�ײZ�Ī6�=�Ϝw;r�u�2�԰��	ix(�ݷK��>    h%ժk�tz�uv�U*ǽ"�kmw�����f���޹G?��߉{-    �� \��W.n:|�����tO�kY� B-tw7�̺��q9��h�3i�i۰�c�����     4�B�u�b4���%W����8֢<�E큳� ����Zڿ���=5�gq�   @�` �����?}m�之�q�e��4�\�R�ujT:t<��t܋B+蕶m1m6�I<   ��5=�:s�u��4>ų��FV+pw��i� �F��+��w��3����^   ��B� 7����U�ۧ�=}.�#�;���d������1��QWƽ0�����u�i۰ix��Lr�   �8����i�k�kv.��9��F�Mk'l�5�q�<����ԣ]�^   ��C� 712��������d�7�=&�;��P��>��:z*�-��^Z]"!����[L=].   `=K����1��1W����|n�J7s���:غ�8�㧺w��k���   �9Qp �2�������>�Mx�I���\��.�]���������XݝҶaӶͦ�%3�    �Z�g��}tL�<�r�b�ȭ�� �~�.����zwǽ    ͍b ��c�O��CG;��.��hZ.���Eױ��Tw���%������}۰�Nq(   �[Q��.�K�\���LmXm�)�]A D� �.L�];���s��{-    �� ܂�??�k�=��j��r'p�����~�Lta�R�{ahA m�`ںIں����a    �gn�5z�u�tካ�cw��W�Lk��ȵ���������x�k   �(3 �=�ҥ��w���R�9�C	���\�b�u��t�x����v��!m�dں�4�QJ&9�   hO�S�G/��g�^�ǵ�z�Q; ��d`~�����3}?�Z    �J ��~��?~�p�o�A"w ��]r7�O���t�8�Tw�?3i�i۰4<d�x�   ���������EW���О��=0�1� b�J�߿����?��l�k   �Z(/ �6}����ɞ?�[H��^���hy�Lu?|<�S��\V�2d�6l��)�    �[�Mi���$�O#^f� b�M{x���?��'�+�    h=� �_���}u��'��q��F���\�Lu?�T�^�UHC�����-�M�=�    4���h:��K��+�*Ϙ�����=$E[@ �ue��{K��sO��~�k   К�+ `�|��C�;^O�Ž��!pЖj�{�,����t&�!vٌ�y�ix(��;r�   4�J�u�4:�:w�5�����������M �Qog�x�]�G>�޿�{-    ZE ��W_=�y��Б����^˵��;��6>%}�M�����1twJ�CQ�e��Jr�   �^\�S��%�XmJ{ƽ& b�,p7~��� �dCin�Ż<��\�k   ��(( `���x0N�ՑS���_'p����r}�ۍs�%Ҧ��ҖM��^��k    V�ܼk�r=jwKq�x+�(j�w~8�� �`������}������   ��QL �*{ⳓ���G�^G�; ,:v����	��q5+��6o\��ޙ�P   ��K�K�����W��I
_NԾ[: ���ؒ?�%�{�ȈU�^   ��@% k��'����R���g	�`Q=p�sW��w�Tw�4<d���N�5   ୪Uץqi�k�41�r2`4�[��~=|e�:13�۵���:����   ��PE �y楉'_;���Bɂ8�A� ��ܗ"vG�0��LC���`4�=���   h7���v�Ҹ�Z�{U���I�����!p�u���ޗ��W>��Sq�   @��� �5��'���c��^�'q��� �,p_��3�͠�I�MC�D��   hEs��Q�~���T�{E�͙$�i� Xc�����)<�§�^�{-    �� ��g_9��#�{�95�����'p�E���\��R�Tw4�dRڴa1x��x�   4��9ץ+��eׅˮ|!���$YmR�*Lk�w XC�a��=�w�ɞߋ{-    �� ��_���𙎃������M� �n5p_�}q�;�L2ii�FӦҦ������   @c��s]�"]��xٵ@Ў&bMj_��})w X#=��]w�>��_�{-    �U �����R�9u硓��]�y�K� �V�/�Q���T4�TJ��_��>d�xh   �cn�ui\�4�:�5����[c&�i��- X�C���[���G���^    P1 �:{���?9x,���ځ'p�E��׹$���Z�Y-އM�� ��   XK��s]��hB�ڴ� �%��j�@�����=��^
    �Q- @>����z�h�?�T��~�� �vྔ{t��\4�dR�8@�   ���y��e��ׅ+�hn�I��<��z�`�����,��/��oŽ    X*�-( hSO�8��׏u�X(ٚι!p�Ek�/Uݝ˭h�T�H�6���D�S   �Z���h:��q��W�����1[�;. �
R	���,��O�~,�    ��k;
 �́W'~������� �V�w X�^��R�KW^�2̤�>��`�o�(eҜj   ��T���(h�<�,��^�r&�R?��, �B�LX}p���}��Z    �zwk
 �ĳ����S}ߜ�Id������8�:��dw�a�r�;kS�7D�{o7�   h=����dmB�i|�U�ƽ*`u��)��[�cg V��+,�ٙ���?5�͸�    7��[T �^��D���C�.d6���&p�Eq�K]�ݝ�g����4�o�8(��$~  ����K���%ץq��l�Xh%�y�D�K� �iC_iv���#�8p&�    ��4�v ���&��o9�{p5{Gw X�(��RQ�.9�;ZX2)���6D��7H�4_�   h9�Ҹt�����Bܫֆ�+h��})w ��7��m��]{F�R�k   �wҼ[W Т�|~�߼y,���pu�	�`Q#�K��]�I=��Ѐic-x��x�
  ���/�.OH�'\W&��IW�����s5j�
yx�� �:2Iw�,��מ�}�k   �� ���K��~�h%V���`Q��KE��ɹd�6�JI�=�Sއ�t�S   �\�&g����Ii|�55����g&��<��F�-�eJ&���)�����~4�    ��h�-- h������ޡ�?;�V�y�`Q3�K���ES݇ML��  �e�����_����OL���{(ܖ�ڗb� �!���;~��O�{-    p�Z{{ ���>���o&�sy2�u���� 5k�T���M%��@�i�_�^�vs�  ��*�Ĵ41�4.]����^���$3W�>���w��Y-޵��c�?���q�    nG�lu@�z�գ�7�6�yr4��v�	�`Q+�u.��Z��b�ud��ӆ~i�@�����   ��0tM�H�S�t�+����`��6�ڗ� nbhCirǶ���p.�    ��j�m/ hB�?7�'�w|�o��; ��    IDAT,j��})�z�N�HRw�44���I�6�>   ���kfN��Ƨ\�є�J5��1�,���q/&^l ��X�]��G�偞�q/    V���� ��<����$��RŖ}�M� �Z5p_jq�������DB�5�I����>��[
��  ��c��)W�������I�����W�0��Ʉ��=��}��ޏƽ    Xl�@�����~�`�W
� ���'p�E��/��3��VH=]�`��  �[�����']SҥqW�����A����� �%�Y�޿�������^    ��� �	��+���ޑ��Lw������vܗ"v�Y"!��D�{=|g�;  ���ͻ&����d�+�����D1{-j�{1��� ���v�Q��>���7�^    �&�� �I}�����9s���춛ݛ���vܗr�����;�G�}�`���W��	N�   �
C���49%MLG��'�\�r�+W=j�gjo�  i�P����V�~������    �-�  ���������M���c��:WA  �su\£��k�ݹ<�M�M�2)�d�Mb&uuH}K���R6��  h�J�O�H���S�J5���� �R&i���k��|��q�    �
�g �>����=�}�X����1� 1�������mˤ��n�`�4����x�  �Y�욚����(h����[@Ծ�жRI�}{����}�}�k   ���V ���N��wf���|"���� ����ָK!�;�"���_����k���z�d��3  �X��53�(f�vMNK�S��B�+�����8�_�T hK�L������=�/�~#�    �Zc[ Z�/����o�Q}m�J��������:�� ��}%��=��`�:�Ro���'���[��t  � _���O�FS٧f��W��ʀ�FԾn����������?��'^�{-    ��b�32���p�����=��:s҇N����|  p_������K��1�vK����n��S��;  ���kv^���Ƨ��}r�U(ƽ2�uԃv��uE���l*]�kca�'>�q6�    �za� Zԓ&��c��V�f����C�vm�2��F�����;�`�d�Ro4�G��^Ϥ��  �j蚞Q�ϸ������W�S-h��#w m!��]�?��g{>�Z    `��� -�ٗ�?��ю�� !I{w���P q��M���z��n\i�A=|���{��.S���p� @��T\�s���4=���Y��\t.`m�$cR{#�@�K%C�gO�_x�喝�    q` Z�s_���7�u���L"'I�6�y�L�c ��C྾�z��eg`]�SRw���[���z�׻:%�  h��kv^�T�Y�ܼ4U�9�և�Ԣv4�	����Ji߮�w�ɞߋ{-    �� �|�KgsG��|��hv�$u�?�P� ��=>��;�x�RRo���G��&��tI�]R"�{ �8��]3�����\�z��ʀv䵨�)�M��@��<X�ض����'6��{-    '�� ��|��Կ;x,�㕪,��~(Ю�\��>��{�f\��Y4ݽ��j����,��  �T�ꚙS��ӳ����\�{u@{3IV���.iSa;@�1I�v����H���^    4�� ��<���񵣝_���$��iz߻�qL ������]&��4�pR��I�}�RO��x)��� ��0t��/�ؗ���W`�(fw�$FM� -%���޽������ƽ    hl�@z�ų�����+��.I�`���e2 �6���.���� [&-uu��;�	�}ݦޞ(~O%� ��|�55#�-H��Q�>5㚞?�	403)�MjGK�@�����Y���?���q�    	[y Ц^}�h���>~����#'}���86 h]�ͅ�h^����i��z:�����N)��{ и��5���检}v�T��y�Z�{� ��Mi7�,9t��_@K�:T�x�����*�    @��2 ���^��7o��d�j�HH�W��;�e�5�7/W���1�&��Ԃ��������RGN2NE k�P�b��S�g祹�(n�|hNfQ�p:����Ԓ�������+����q�    �|  =���y�hׯ�僤$��iz߻�q� �Z�[G�K!�݁�RgN�eM�(���4uu�j�V ����k!_�֯��g�\�r�+�*L
T���)b�!pд�ٰz����?�T�W�^    42��  �����廾���_\�LwK��Ӈ�(��X�u���z��b�;���Z��a���Rg���#
�N]�T���i~A��K����Ř=_`
;Ъ̤�����hJ��s�l+>��S�ߍ{-    ��� \��G3/n��ɳٽ.WGN���	�q� �����tw��<@{I$����'�wv�w�D�; ht��kv^��[}�B^�����hLi��q �\\ڳ�xx(�}�ȈU�^    4� o�ԁ��8x"��Je�DBz��@��s		@�#po?�dwɝ�� �ͤ\fq�{GGm
|Δ�FS�s��c^, ��j�5��b�h�צ��&��j5�U�S����pc<��4R	�ݻ���������    ̈́�A �u}�KW~������|"-I�w�~(Pp� мܱ8ݝ��~l�L&���S�夎�զ�KݝR*�y1 \�Tv�Q�>� -�������ϻ�E���S�q�8� h
]�j���?��'7�N�k   �f�V! ��^�����Ѿ�=��*��{Mz��N� ��;�U�݉��v���}9�)�#M�f��)��:�V�㥎��Q -�\������B������_�{Ω ,W}B;A;nG ohCir�����<>|*�    @3b� ���xn�?>��+UY*)���ڱ��O ��;n&��%�q�hI��/W*��ٌ�#'ek���>��2i�h ��jU�P�
��P�"�B^�ˢT(D�+����ip �3�ILi�j�a;��efڽ��گ>��`�k   �f�6" `Y�������B�$$i�N���Ȍc	��A��[�^���!��}�� 
ݳi)�5e2Q���>�V���-��<��U��|>���E)_\��BI��]���h�V�X&�9A;�JC��h_���{�\x��O�?�Z    �ٱ� X��������ܟ_O�J�`������x�9��vy헰�hF��ߪD"�߳�(�Ϧ�L��[����NG�NK?�
4�rE^,IŢT,G/%W�$
R�T�y�}R�槺��13W@Ў��R�� ZC_o�߻��w���?ǽ    hl3 n�Ȉ���֑�����ʤ��@��M\���ܱZܣ���&�:�$Z+p��d�G7[|=�]�3��m�a<�R劼\�JKnŒT,Gaz�M\��������o�;�E�tv�������4t��S��=�c�mY�{9    �*�r ܖO�t�ŃG;?^(��tϾ@�c� ��kŽ~3�����v%R:U��ҩ(|O��t&z�JJ�T��?6��>.��1�ۍ�R�U*K�T*�n����%�Z܁v����H�'�� 4�TR���o��L��Ľ    h5\�  ܶ~y��?���L*'I�6�~�}���/ �;փ�~	k�;��FA��t*� �LH�Z$�LDoK%�P~���L��S	)��&�[}l"�Ty�X��j5���U�Z��e�Z�JW�"Ujo���W�D�>�U�H�j�>,E��3�T���Gc��@�z{���w�~��'��0�    @+bK �"���w�����>���re3��7�M9� h<����]LxbD��jҩ(�K�� !%�TR
��ۂ(�OԢ�T2���cLA����jD6���/�L&$#�_�zd.Ia��u�Z0^�D�+W����X��UKe�C�\�����T�\�*U��j5
ӫa����܁���A;G| �qi���w�1���۲�r    �U�E	 XO�4�k����Ų3�����or�5 �;E}��ӈ�����/���fє�����Z���������{�������<�<�r��_W���hu�� ����$cM�s{ �H%�w���뗟����    ���J ���ܫW��G:���L"'I[7�>��R)�7 �;��	���Z"p���dhnLhG���������S��g���ø�    �-L ���җ��\���S�ٻ\RgNz��	�s�?w4��J���m�.�� p��#p�I��	�т8��~,��M�s��]���G���^    ��4 k�S/L���;~�X� ���}_��vs)@��ь���w X9NF��fRP���.Z�� �E:�ow�_|��Ѹ�    �-N ��y�+�y�D��O%;$i�6��J&9� ��;Z�;p��`�8� 
A;��� �\ow�p�so䩡?�{-    Ў�� ��/}�l��D�_�8���M��I?���6p���ъ���ׂw��7B� +G���$��"p��,��M�s��]���G���^    �+�@ ���&~�����I����~�8XG�hN�\�; ��;��̼�������H'�������?�Z    �ݱ%
 X7���#o�����D�$m�h��{e3� �w�����LN��E� +G��%3�Ąv`8���z�*�{w�����m�k    � ���/_�<>���S��}.)��>���l���G�D��}1|�!��; ��;�jj1{`������t���S{�~�g�^     )  �<0������J�Iw�	��{MA��	��!p��k�D��Q
�E��������������H'C߿���_~���^    ��F ���W/�w�t�9%�/I}�G�������A�,_}���jSށfG� +G�,�b�n�,9.�����b=��={�?���}�9�     ގ �X��x0L�ё�G*�,���/�]��e`���/���wr4w X9w�z���;���63i���kC���#�Z)��     ���V @C���㏾y"�k��$��j��wJ&9VX=���b�;��; ��; ��s{ ��+땻�,<��'^�{-    ��c� �0F^9����ο<}>{�$uuH|_B�9^X�����/Q�nh0� �r�h?KcvU���=�[�y�4�kg��#�8p&�     �{� �����&���';�Q���L�������"p�_4�����9�C� +G���Mcw��� �� �-�t߻���~����Z     ���, �!����?�����JuH��F��(���������S�er��w X9w��$�ڄvbv��pn`Y�{*�{w���'��0�     n[� ����G3��7~�ȩ��Bwe3��hx��w�q�c������Y��L�Z��W2��8�pS&i�����~`�^+Ž    ��c ��}���^?��ɅB�0������MA�q��!p���~!z��!p��#pGs����-�s{ 7ԙ	+�w�}�S}/Ž    ��ck �>��.�>v0����!���c��{��p,�|�@s�G�D�=� �r�h<��@[���um,M��1�#���{-    ��a� �T�<0�?>���bEA"!=pw�����c�e pZ�բw&�cY�`��'��]��elm�s{ o�J��#�_��o�^    `u�� h:�}��G�����NI4}�uvp\ps�@{��/D�x+w X9w��$s��dv �ù=�������v���sO��~�k    ��� Midă�`���~(�)���s�=wp���������xH�n�`�ܱ���쵉��� X���̴s[��C;����c[�^    `u�U hjϾ2�3��w|mf>HKҎ���
�Nq��v� ���K�QI�4w X9w�L��Ո���m��hsٴ��w^~��}��{-    ����1 ���������>;�����e�|w��M\&�V� ޑ�c�����^V�; ��;��ef�1�q1����hc��J���Q��g��x�k    ��� -��&�����/��0������; w +�8�]��̈́� V��o����� ���@J'C߿���/?��Ѹ�    X{�5 Z�s/��{�r����\�ݦ�7P/�< � V_}�;�ޛ�; ��{;��'����@,8���Pizǖ�=����Z     �-h @Kz⹩�?|2�_W�ff���=��$�}@[#p�^��K$�#p��#po�����ޝG�y����w��>ҙ�Q�lK��Ĥ@Ka5we��i���6-�I ĖE����r��1$���қ�B�%�����;	��dk������rd�vdkK����|ֲ�s$Y�d����~��){�f�p+;P�d{(��r��Y1�����  ��+�{  ����o���?��?�e�w��G�g�Z~  W^���'M#Ji�4�r)�Rz����Ҙ� ��$"��|.)�Y�J��R�4"}.ψ+ @z����qݩRn  (&�M��&'��Trꏾ���}����#�)����E�PDnp�����/���<<��w����F�Fv�	����J�$[56���r�&'����   ^��6~�ďm���'N��cCI���4����P$
�@��Pt�P��,��x��.��{=��"{����	��Ф��g֯����_���g   _^��0>�ѭ����W_��E�U#�p[�CֽP
�@SH�+�?_z����~	�.��{�+�'�=_^��P@�=4�$�X51���o����l��   �?/}P8�>�3�쒏�:�V""��%q�iTZ<��)�Ep������<
� �O��jH"{�����ؕ�^@��&ұtav��ٷ���ݿ��,   �/�PH[�X��t�K��\r�b�E[5��[��2�f���E��G\(�����p��k)��H�ؽ*pId{hI�Ĳ��[����s"�y   �/^.��6>x�޿�^���T��6whv
� //�.��~��Y��F�.����u�6����#��j@���^]�[�r���ջ9�Y   �O^J��&�����/m�]]�%�6whb
� �^vQud1�����]���)����[�#���^Q ��d{hTY������%go��>��8   �//��s6>xl�S϶����6whF
� ���[��[�� ��p�
Zp��~�6v%v�: �C�V�[1���ݻ!�Y   �^�����ѽ{��~Ǟ�J��C�Qp��^����%�<(�\��-�'�;@��$i�L\�l�6������  �1x� ^��Ol��g+�85]r�;4w��r���ϗ៻���._�ܳH�$.<a..�+�4$�D��-�[9��n����g  ��x� ^�����}q���Z��CsPph,��/���b��_:w��W���O^|��@3���]��}b�nz{�ּ�  ��x} ��w��o<۶��T��6whd
� ����>y���;��ˡ��|I�E��+��lu�Z]\�fb�׶l�}[޳   и�  �L>���౥_ھ�mm��ܡA)����{�e������_���# �����7�?�G�ܼ��Sp�:�$I,�ڱ��?��-��  ��fO  ��Ƈ���϶N�>Wv�;4 w��z��s���e�;��.���E�\C=����Ba]q��Pp�:�^]�[�z�}n�yo޳   �� �U����݇��ǟݽd�bns���PX5)�|��������/�{�hJ�ߴ�\��?��u ��u"��e#�;�[�y�;~&9��<  �S�    IDAT 4; x���Љ��ƎʇN�)U""V-K⎛���L����j�[��qq���o��@��ԟ�������|� o
�P:�.�\�b�޻���y�  @� ����~�p��v�m�n1ˢR����4V/w�;�#w�ª��+��]���	|;߼Y����9���\އ� �[]�{hv�4�VML}��w~����l��   М,# �����}z[�G��J�cCI�ykK�<k��(�VS`^����_����E��E�������+� ��T�IW���u�f~��=��{   ��e ��cYV���O��7v�~��|��K7�K���W�<)�V�0/Uv����/�3����� ��E%���Wz��/|�����B �]��=\m-�$[�|���h����d>�y   h~� Pc��|㳻�;x��3"��;�7ܚFO��.�M���`.��2�K�_��Eo|��$�o�Cݻ�{��r��~���F�,^TFo�rz-�g	@=���*��^8�zb��￻�y�  @qXF �����~��g��if.I�$���iܺ>�R����PX
0u��n�qY�%�|�/|�h]L/,�G��x��_�H^�wKa���W����p���5�g�������y�  @�XF ��GO�۶#��][G#":�F|ǭ���<(��LA�/����|����o~��~��$��/E�����ɼ�/Ћ�����%~���3����.*���/e1�� @��{��{fO.=���7�E޳   PL� p��������35���$b�DwܔF�ų�&w��R��n���|�K������p� �� ț|WH����v��o?����,   �e \%���О��/l�Ӷ6�,ڪ�ݐ��	��Z�
K�v�aț|5�$I���]>�����޵5�y   �2 ���<t�����Щ��ֈ���$��4��<��JSp(,��qv o�=�P����k��>��ޮ��   .�� �<�X����O?�}w����K7�K���I��3\1
� �� P;ά �M��(��l���_��X��L^���=   \�2 rtߖ#?�coۧ+wFD�&������W��;@a)� Ԏ�* y���2�uϝY3�������ټg  ��b u�������wV���LRJӈ�M��k�HS�j�%w��R���T �&��k�V]\X�|淶l���y�   ��2 ��{>�{����۵�myYt,�x��i�%��P#
� �� P;Ψ �M��W)����ٽ�#g�{�Fv�=   |;� Pg6}��۞޶�'ΖZ#"�G����4��<��r)��@�8��7�^��+��y��ޏ�=   \*� �C�<��mש�?޺�����Hʥ��פq�I$��7�V
� �� P;Τ �M��K�Rʲc3_����>��{   x5,# �����c�������w��IDOWwޒF�g8�
� �� P;Σ �M��W��1�;}l�������/�=   �� � �y߉�uW�[�M��$�X9���7��Z�,�WC���` j�9�����2�Z�[1�n����g  ��a �O�{���/�<P]��ET*7�K��UI�g:\w��R���O �&�Ë�I��g�Z�����g�cy�   ��2 ��G��Ķg[���rGDD_wwޚFo��:|;
� �� P;Ξ �M���tw,L]�b�m����ɼg  �Z�� �49������mW��g�4I"�,O���(�=���(��@�8s�7�"��%[\=1������g  �Z�� �����^{h��v�.�"��q�i��H"�o��PX
0 ��	@��{
-I���;8p���{�o�   �� h���w����#�O��""������4:�=��b
� �� P;Ι �M����;�VOL���{�>��,   p%YF @�����S��۶��g�4M#�Y�ƭ�(�<�!B���` j������NkK��j���~��v�1�Y   �j�� �&����ݶ��s��U�gѾ4��7�1:�x�Sx
� �� P;Ζ �M��0��blxn��������g�   �� hR�y���m�Yy���R[D��@��%��v��K���` jǙ����B_�ܙ��f�����O�=   \m� ��&'��Tz����\�3s��i�5�Ҹe]�@�(��@�8K�7���V�..�Z6������   �b ��GO�۶{�w�.�"��q��4�,O"�(w��R��gH �&�Ӕ�i�-���5+���;~&9��<   �'� (��9�Ϸ�j���c�Έ���$^wK�=2Š�PX
0 ���@��{�N_�ܙuk�~z�[{�[޳   @=�� �����uG�O��N�I�r"��oH��U6��)��@�87�7�����uq~�����{��M޳   @=�� ����'����wꏶ�n}��|����צq�5I���@sRp(,��q^ o�=�\ʲ�c3_����N�=   �� (��9��v�o���[#":ۓ��$F�9����PX
0 ��@��{W��p���ё������~1�q   �^YF  ��۸mg�='ϔZ#"F�x�-it��4w��R��gD �&�Ӑ:�.�^�l������g  �zg <��ں���g��]����$MӈkV�q˺$�e��Ƨ�PX
0 ��l@��{J�������|��v|����l��   @#��  ��;u͎}���{+��$ڪ��Oc��$2����PX
0 ��L@��{BY���8���=�7y�   ��2 xY�=r�-��(�ȉ���,���x�-i���4&w��R���A �&�Sߒ4���������_��L��   @#��  ������7vV~��ٴ%I"V-K���hm�%h,
� �� P;΁ �M��nu,]�]5>�ч6vߓ�,   ��,# �K��#�������m���;3i�q��4n�&�rY��1(��@�8��7���S�,.�������&'����  �Fg �*}����Z�`׾���H��Eܼ.��˓ق:��PX
0 ���@��{�F9M���魫֤�s�[��=   4� �5y�O��g�����?"��#�;nLbd(�/�[
� �� P;�| �M�'Y�p�챉�����{>��8   �l,# ��r�����g�V7�<�V#"F���4�:�ꏂ;@a)� Ԏ� y���UO��Ԛ���y�;�>��,   Ь,# ��69��g[N���;�?:5���$b��$nY�Fk��A�Pp(,��q� o�=�Xں8�z���l���Sy�   ��2 ��Ϳ~ph��?ر�r��|����צq�5I���A��
K�v�� ț|�U�Rβ�3_����N�=   �e Ps����xמ��{�fIĒ���ץ�fy��A��
K�v�� ț|�U�$ˆ�w�����;��>�y   �H,# �+f�G~z�����Dd�ם��7�1�'��w��R���9 �&�s��uϝY�l������t޳   @YF  WܦOl����_8y:m��H⎛���E���
K�v�� ț|�ӱtav���Ƕl�|g޳   @�YF  W�cYV������3�[`j&)�i��eI�r}����C���` j�������\[���ʉ��v-v����d>�y   ��,# ����ǲ�mw��޶���ΥI�%��k�X�:�4�M���
K�v�� ț|Oʹ�#[6:�7���drr�P��    �YF  �x�ߝ�n����w��_��}i�-��X9�D&�p�(��@�8��7���VN�llhj��h�o��޵5�y   ���  r�+<�}{T>��`�h]Iܼ>�e���B�)��@�8��7���,�,F���������|��    /�2 ��}��]�>[~���JGD�I�zC�}�
���PX
0 ��@��{^�,b�w�䲉������O�=   ��,# ���a�_}fw�_�>W�DD�$q�Mitw�-\>w��R��g3 �&���uϝY1:��{�>��,   ����  ���d��m9����Yy���R9I"��&q�i,]"���)��@�8��7��K�վ8�|d�׷l�}[޳    ��e P�&=�~�H�g��|��l��i��eIܲ>��V9�WO���` j�Y����������+��|�c��͓��|��    ��e P�6��������`瞖�f�Ӥ\��vu7^�D�,�p��
K�v�� ț|�K�V���i�m��n�0p:�y   ���2 h����v�+���=��#i�D��&�u��HS��oO���` j�������@K9�e����;���ѿ7�y   ��g 4��?|��=��>��@��,��m7�Kc��$B��(��@�8s�7����(��l|pj窡����_�{   �v,# ���qˑ>x��k{�g�Ց���X6��8�$w��R���- �&�]1�?{l���OlzG���   �=� ��m�r�v�i�|�xkGD��I�vC�}�/��PX
0 ��@�����"f��Y�����?��8   ��c 4�{7{ߎ��x�dyID��H7�K��K��<w��R���+ �&�M��P������M������   �<� ���}�޿�`�[/�G���FEw�
L�v�� ț|_ =�S+�gx�]���   �z,# ��u��O~����N�)�&I��p��O��S**w��R���) �&�@O�����l�����g   �>� ��k��>���gO�)�&IĲ��E��vY�h�
K�v�� ț|�ĺ��Ϭ��ă�~1�Y   ��XF  �09��S����mg�'�L�Z.�o�>���2QQ(��@�8?�7��	u-��Y>1��-�����g   �g �cYVz򁓿���ʛ�N��i�b<���St/w��R���& �&�7�Υ3+��w��Ο�{   �~XF  ��eˁ�����=����S�i�B���ui,]"#5+w��R���% �&�7���ř�cs��   �K��  
�;�|b۩?ع�����(�i��eIܼ>�j���l�
K�v�� ț|��:�.ή���[6�(�   /�2  "},k��N}晽�<=�R)bՄ�{�Qp(,��q> o�}j�.έ���]o��L��   �o�  y�����o���gw��qj:-��kV�q�5I�*�7<w��R���" �&�7��j6?16��u��~䮻F��=   �,#  ^�o�v���֓��c�wM?Wt�vu7�M��E�jT
� �� P;�C �M�o K���?�zS�L^���=   �X,#  ^�䣇�O��Ύ]�rv&)WZ"�]�ƺ�IT���;@a)� Ԏs y���X{uqnbl��G�soڰa�t��    ��2 �L>z���і��cO����.���5+Ҹ�$��2U�Pp(,��q� o�}j�.�M������s?r�]���   hl�  ���RĪ�$nZ�F[U��w
� �� P;�= �M��#�ms+�g�G�Bכ''����   ��e �k��/g-[���޾��#g��r�F�O���h_*c�+w��R��� �&�ׁ���3��~w��Ο�{   ��XF  \��O�[r�`����[}㙩��B���k��h��ꍂ;@a)� Ԏs y��s��=vbh����}O޳    ��2 �˲�W8����V�ęRk�D�'q�4z�d�z��PX
0 ��|@����-I��k�̲��?��羼�   ��e @�ݳ��C�����ʒ$�bl8���K��[�ʛ�;@a)� Ԏs y�ﯖ,��g�̲��<����y�   �e ������C�o?|��3"bd ���O��Gˋ�;@a)� Ԏ� y�ﯴ,b�w���x�{7t|<�q   �ⱌ  ������_ڽ�������,��K�k�Jd��L���` j�9����WHY��[><���o��T��    �e p�l�����@���f��ǆ��䲫B���` j������5�D���������l����=   �e �Uvߖ�?t�p�c{-_X\L�z���$Ƈݯ4w��R��g �&��H��������z�;�?��<    XF  ��=�}��C-�~��։��H:�F\�&��+�HS9�JPp(,��qV o��e���llpz��p�S��bדy�   �b�  9����k����]�[o��KҶj�ڕi�_�D�,�Ւ�;@a)� Ԏ3
 y��_�j���������4���]y�   �r,#  ���ç�O�]��v�~ϙ��R�X�"���&�V��jA���` j�������R{�����쟏T�޴a����   �v,#  ����f�����'w�-��ԙR%M#V�'q�it��o�C���` jǙ������k������ݲ���   �հ�  �c�l>�О�����J{�d16|����#ǽ
� �� P;�" �M�%YD_�ܙ��o������   x-,#  ��|��/?{����G*�Y1ؗ��&16�D&�]2w��R��� �&߿�r�d#�3��O̿u�[{�[��    \� �r߇��y߾�#�WF"��Jb��$VN$�ݷ��PX
0 ���@�������񑹭���?y�ۻ���<    �` Ѐ6=t�<^��}ZW�-$I���uk�X�<�RI�{9
� �� P;� �M���%�labt��/O~잷��{   �Z��  h`|��Ğ#-�ڹ���N���JĚ�i�[�D�U�{1w��R��� �V�|߱tqv|x�����]w���{   �+�2 �	|��Y˳�;���Z~�ĩ��r)��+�X�&��Kd��
���s�  o���I=�S��ٲ���   �J��  h2<q��#�;j�$bl8�u�����
�x�+���
 rW�|�F�}s�FF�&���cy�   p�XF  4���g{V��26�Iow��$�b<�$)fTp(��` ��B�% �+M��+�,��>1����wt.�y    �6� �&7����=U�Ԯ��wLO'��j�ڕi�[�DKK��;@a5}�**���Դ�~I5[��Z��&�޻+�y    �b P�>��o��ص���N�I[�刕�I�[�Fg{1r��;@a5m �8; Pך+�g=��S��Y:����d>�    �f P@�z�ɏ�>�����*I1ܟĺ�I�%�5qFTp(��*� �i� 4�����4Ɇ����/l�Cϧ�   ��XF  �����N�>��@e��|��t%q��$VN$��͗�
�)
0 u���	 4������lqthv����O�����=   @=��   >�[S�vl���;�U���TRn�F�Z�ƺ�IT[�'3*�VC` �LӜ hX��;�.̎�~a�:��N�=   @=��  �y�eY�8�]���ȉJG��|,��I���񳣂;@a5d�N5�� ���0�>�,�{�N��,~���vm�{   �Fa �K���#����_�{�:>��`_7\���PY��Hw��j�@hȳ  M���}Ky1��9�o�����=   @���  �=����w�_����;���RWG��&�r"�4m�<��PXu_�h u �)�m�oo[�����Ι������y�   Ш,#  �$����:���Ww�/�豓�%��,��%�nm�퍑+�
�n0 �!�? M���}��9?51��so��L��	   ��YF  ������m}���-�YD�'�vU�F��:Θ
� �U_��V�y�¨�|�RJ�ၙ�C�s6����y�   �L,#  x�����;�/~r���S3i�ciĚ�i�]�D������;@a�E�I�]��pr����k    IDAT��l~dp�������u?��,    ��2 ����/g-���ɏ�>X���'[;�4��cI�_�Fwg�dNw��Rp����� �U��ID�̞\�/n������   �e  5�iˡ=x��y߁�Us��u'qͪ$V�'I���l
� ���P;^S oW-߷UF�������������   �e  W��C��O�T>�ko��N�+Uڪ��Z�ĵ+�X�$���
K��v��@ޮl��"z:�Ɔ�>w�๟���sW��   �[XF  pŽ���>p����w�b���p׭Jbx ���T����j�k� ������b6:0�s�g������ؕ�1    �4�  ��u���������'�;����g�׮Lc��$ʒ)    WYw�������u.N�err�P��    �� �UT��x���hG��3v\_�zG|��X1�ĵ����t!$    WN��P�졡��������   �Rp �K�,�ˏ�c�ǵc�q���ٽ�mg)��X�"��$�4�I   hK���#��7�9�/6����   �)� ������5�:�qj��c��U��'�D��jYk���ў��    4�4���;96��_�s]o��L��	   �W�� @]Hb>��7O�Y�M��='�{㩭Y�'�fenu   ���d�ó�ӿ����R���=    �N� �������gbew%N�~wl߷2rIT[��   �KJ"��c~jlx�s����ްa�t�3   ��)� P�f���'q늈�ŵ������~��   �%�ladp�ޮ�������=    �G� ��PI���ޭ���-��|O��?_|�mnu   (�4�b�o��`_��-;ߙ�<    Ԏ�;  %M�����ѿ2b.[�O�۶���>]���$֮Lb�D�Rޓ   PkK����_���~��ɼ�   ��� hX-ɳ�����L���wƎ�k㉿j���m���$�]�Dwg���    \���b������G[���{�;����g   ��Qp ��I���ㆱ�㺱�8t�;b���غ���[�   h]�|x_���i���y�   �U�� @S)Ǿm�L�^�Ĺ��b�����_w�מJ��]�   ��]��}E�W���m��    �w  �S�Œ�W����ڡ�8t�;c��ш��=    I"��s*V�쌞�#��G    G
�  4�$;CK�{���Z�-vY�w��B��h    �U�,����1��d��;ο3�u$    ꀂ;  �Җ~5��j�ZG�}w�9�,��ڝ   \i��P�٘�-�GY�b�S   PO� (�$;�m�3�'"旍ǡӯ�]������   Pk]�11x(��R�{    ��  �W���h��]1�xK�=v}�=��siޣ   4���B���ޯDkl�{    ��;  \�-�Z���Z��o���� v^����b��=   @�+�Y���C[cI�x��    �URp ����TtW�$��"�������Ǯ�CqzJ�   �X]3�lh��y�⩼G   ��i�  ��Q���h��Y1��.v�.W�   �ձd.&��P�_F9�}�����   @�Sp �K�$K�'��'����89wg�=�2m��[   � ZJ�1:p*F���'ο3�w&    ���;  �ILEw��{��~�7�L�!v��g�"�lu  ��&}=�b����~1"��{$    ���;  \�$��@�gc`e�l�"���-v���S�6   и��gcb�P�)�q��;��~    �0�  ��J�#F�w�Ț����b���c�Θ�O�   �۪Vbb�H��|-*��y�   @)� ��$m��ƚ��ƚ�R��C�>�&��ż�   ��J9���31ѿ-���G���   �#w  �����x�~<֍vǡ��{�Ʊ�U�7   ��J)b��T��=�忈$��{$    �w  ��O�`�gcpy�b:�N����3��2uw   ��I�,���b�_t�~!J�ټG   �o��  9I���ߏ��ي8z���}p0N���=   �$���ꘉeC�c`�#�y�    �H�  �@%�#�;b�=b&[O���Ź�Rޣ   �B�}|�pv��Q��=    \2w  �3��S���X�1�����b��ޘ�Uv   ^^{�\����/GK<s��Y�3   ����  u�OŊ�bYwg^������cv>�{4   �����������$O�=    \6w  h id�Qz":������8�����8x�=����   ��j�B������y�    5��  &���*�Yt�D�i���o�}G����K��  �I��,�����y:ڒ'#���   Ф� ��%1ݕ?����qj���{dU<�s��   ���*1�{:{vGW��H���G   �+N�  �E6��/D����89wg�?�B�   H��#�'c�gk,-=idy�    W��;  4�$������=��   P��Zc����R{�D�i�   @~� ��)�  @�YR����S1Գ5:JO�=    �w  (�o)��G�?�,m��9��  ��Աt.����P�_G%����   ����  ��Tt��,�#������q�����+��Jy�   M��m.���p�_E%y:�q    ��)�  ��'����X3����q����{�/�L)�  ��J"��}6��N�p�W��l�{$    h(
�  �eYT��ǲ��ǲ���XGN]���Ɖ��Y���   PW���ꘉ��1���(g��	    ��;  ����T�w>����8t���w�?N����;   EUJ���>#}����(ǡ�_�    �E�  �d�dk�wn��Έ�lY>wk82�NUc�  �&W)/�P�����-��l�#   @�Qp  ^�R�+����Y�'gn������Θ�O�   jbIu>�zO�p��XZ��H���G   ����  \�$;ݕ?��Jqz��8t|u�?�Sӥ��  �K�DDg�l�����������	    
E�  ����(=�O�����XGO��}Gz��jdY���   ��4����=}K��l�#   @a)�  WT5�����b�#b�4G��{����KbQ�  ��T�Y���ួ�Y�_QJΞ�
gU    ȕ�;  pդ{c�mo�G,Nt�������q�Ē��K�  �&ױd6�{��P��h����Q    ꎂ;  ��4;}�?������$f�����k����8u�5�̕y   \�$"�:fb��X��uT���	    �6� �ܥIm��bY��bYW�|�<���9������B�  �(*���;�]�����H�X�#    ���;  Pw���Z�3��FD�$���OLā��qn�1  �oJ"��}6�OF׳���d��o   ���G�þ��������q��ծIˢd=�� 	���[��}01>I��O9&�!��#�iŴh����(��.�ݙٙ鞞~��aI�E��Hv����a��k���bf�o�xX)C  �v��t��ɕ�SW�U>��習;ws|6�F�   ���Uuw湺7��?O����    ���  x�T���[�>I������գO���q��r��  �(��N/���I��|;�⹷��{�    )w  �U�^��-�ד|�Ȣ�b��r^��g�;  �CΖv    x<	� �GC�dP<���sc�ԙ�|�ky���ܾ;�b��  �6+��L���w?Wv��q�Y[�   �1��   Ieγ����\I������?�W�����8�z�  ��69ܝ�����M����H    ��	� ��B�[yrt+O����(��_�맿�׎v2_��  ��P$ٝ^���q�L��~�KY�qҖv     w  �1Tf���g�J��+�*����/�����=d]�?�&   �'��:W����3��E:9��H    @�	� ��^�������>Nr����K9�=������l��A  ���׭s�;����9=�*/m{$    �!"p  x�M��s�1}.7�ɦ�b��~z3����t�O�(�  ���$��<qx���w��s)�a,    ��  ��b�I�k�$�<H�y2g�����_˫G;Y,U  ��H�3Y����\�y%�Ο�(�    xD�  އn^�~��g���3O$�|*G�����+�{2�jSl{D  ��h��ս�\ݽ����S�h�#    �(�;  �ϡʭ<9��'GIs��l�k9:{*������A�f�  ��^�+{繺�Zv��*?��H    �cB�  �!)�ʤ���i��K��s��b���k��rt6�  ���4�/���I��I?ϥ,�=    �8�  |D�\f��zFӯ��4�3���˹wv#�����Y/zw  `z�d�"������a�/S�m�     p  ���9�N��s�|��A�>_�j^?���Ovsz.x  >ݲ��������2��E���=    �;�  ���y&ݯe�f�^���Ws��Z����l^�i$�  �����9ܛ�p�8���7Sz�    x�  Z�l�e��?��O>}%i���V���Oo��������I��1 ��Uuv��\ݽ���w��s)�mO    ��	�  Z�hN߶�}ӌs��r�f7r�x���A�Z�  ��~U�`g��ݓ썾'h    w  ��D��=�w��v�&U�r4{&�������,7۞  �(��_ݿ��ѭ�¶G    �H�  REV������ܘ&��*ͯ�����;����P�  ��p�Ý����n�T���=    ��B�  ��(�ʨx6�鳹1M�N.�����rt�����,.;�  �1����d�����O^ͤ��t�ڶ�    �
�;  �#k�a�|���s}��Z�.��|��9>����wrz�O�l{N  x���:;�E�������V���m�    �
w  ��H�����v��O$�f�y���_�Ƚ�{�w�����  ��(������r�s7���3�o����h     �$p  x�u�Y��?�t�\�$����.>�{�Wr��8�E/Mc�;  �ݲ��d�����^�n��9��X     �;   oS�V�r8H�D�)��l����]���n����a  �$��:��Yw��3�nzy1e< 
    �A	�  ��:͝�Uw�w���A�t��/g�x:��9:����'� ��W&�N�9�9����L��n^��X     ��;   ��&������[ޯ$��g��B�����N���Y��m
  X�d2^eoz���qv�?Ƞ�f���=    �#M�  �ϭ��L��e��<���ئ�����r����s:륮��
  �_�ٙ.r0=�����V�H��m�    ���  ���d��J��I�$)G�o>��������l��E�fۃ ���Wu���ٟ�fg��L{�J����X     D�  �ǥ�gT|=�����8ɵ$�N�V���ō�����l z �CUu�G��Ogٟe<�~y���    �5�   lO}�i��2�$�'I�%u�2�|�m���E��I x�I��ev��6f��Ŕ
v    ����  �V)s��}S\��곹?{2'�Ӝ��s�*�=*  [T&����ߙgoz�i��/�(��    ����  ���4w�۽�����ǚ�|���6���4��  ��n�d2^fw|���<��3��U�̷=     2�;   �"G���^g/��g��_T�� <<�U���2��E�'G��^^L�:    �ǂ�  �GF��wD�)Y4��������l��Y/�����  ��~Ugg����<;�W3��u���m�    �	�  x�5��B�r8Hr%iRe�|.狛9���t6�鬗����  ��N'��W�Ͳ7>ɴ���;�J����BK�    {w   ;EV��p��\&9|p��A�7����FN�ws6��l^��� �=�v�LF��OgٟeԻ�a�[I���h     <�   ��"G�v�,�Ir}���A�Og�|����l��y߶w ���$��2��";���e�)���w^l3;     ��   ~�f�A�|��s8Hr��𦸖���_<���$g�A�/z�l�:- ����&��:��evG��eX� ��V�/ׅ�     ���   �t�;�Vw2��L�:�in�b�9[\��|���a��}�; �zE��`��h���,;���ng�����o{<     w   �u�W2龒�$�>y�������3�-��t6�ټ��y�M]loX �կ�L���N.2�f�5����w^\��    ���  �ǠS�����Uɍ76�7��l��|y3g�����r�d>�n�;/ �h�6��V�Nf��g:�Q��[I}���     �'�  ��Y�_��~������y��e��\ln�|~���8g�a�U�k���+�d<\f:\f4�ggt�Q�N��S��/��    ��  @�l�+��^�;��I��֙&Y�Oe�����nfÜ���]T�� mU��x����"��EF����A�:�f��    ��B�   �"G�G�����(G�X*����.vs�g>��⢗�� �2W��.3�g<<ͨ��a�{I}���     �#'p  �GA=ϰ|>���9��ԛ[����/ws:�<��>������ ��~Ug:��xt���"��݌����wS����R�3    �6�  ���[���~?�1}�ܺ��,V73_f���|>�����E'�� >�"ɠ_g4Xf<Xd<\d�?Τ������Xl{D     h%�;   <ƺ�˙t_Τ�d�d���:E6y:�뛙-�3_�3�f~�����զ��� �
U��`��dx��`�q�au�Au'U��Ym{D     x��  �w(Ӥ�K��/=��Go?�� ���,VW3_�fv1�l��b����k�; ���Sg4\g�_f<��h0˸w�~�v:�����    ���   xߊeXe�O��I�o�k�n��ӹ\_�����n�+%  ��-��댆ˌ�����{������f��/�-     >tw   �CU�T���{�'n�4㬛�r�����~..��]3_����r�,�ler E��ΠZg8�d4�Ȱ�Ƞ�a�nzݗ��k��bߐ     �c'p   >V�b�N�b��$�$㷟oR�n�̲����j����.����Y���XV�l�19 mSɠ�N��d�[e<��h0K�:K�s�~�Rʜl{L     �}�   �Rd�N�J��+���~��[��i��̓�\�e���b9�l����b����&��� ?�"I�Wg�_g4XfԿ̠w�a�~��{���?}�:     �P�   �2MR��Q^ɨ����k�:�;׳��e�|���_�U����庳s��.WEuyYv��c�$eQ�Wm����2�/3�/2�f���e�y-��0EV�     ��	�  �GNY&es;��v�����������I�����u��Zw��Y57��'.Wٹ�,��U�w�,��(u� �MY6�W���{����wW��SU����)���NYn{Z     ���   �c�~��O���Ϻ���z�F��.�/o�|�򲸹\��rY�\.��jUV��Ng�i��al��]Q$�^]�{�NUm2�-3�/ӯ��Wg�wN�+�h^���z�D�     ��;   ���o�ŕ&�/o|��?��?=_����4��7������r��պ�.W�x�*��eQ]���jSi�� �U�i�*u�m�U�^V�f��g���W��V��o�����_���|��_�������7��     �s�   |H~��v�������?���^���AV͗֫ⳗ����2W���/7��j�W�n�Z��^��(����)������ͦ���_/���{�漬���6�    IDAT~ռZ�~���[e���t�z�w��ٶ�     �qw   �-�����<��z��=�����߿���X�ͧWu��eqm�.V�fg��L֛b�\wz�U��u�Y.������Qi��JSu�ۮ��u{9�ͽ�jn�����7/�Ο��     �CO�   ��W�l��$Ͼ����<�T��K���ӗ��B�yb�ɕ�:��:�ͺ����eo�)��*�զ��uQ�6v��QE�Nݔ��U��t�f��6ˢj�����v�YU5�e�>�:�kI^�������6��o}�_^�ֶ�     ���   a��O�n%��A^��o6�����j���j]>���yY��&�ͺ3Yo2���p�)��:�z�j��t6u:�Mѩ�)��Z(�C��ISM�ݦ.��e�4U�Yw;�����v�E�S��Ns���)�{���]Ty�����~�7��     ��   ����b���o||��|��V��/����l��̲x")�^�y"�b�n��jS�d���u�_ם^ꦻZ�_7e�٤[�EY�(֛t�MQ�u�u]M�|8o��JQ�u��4MQ4M��M�ɦS4u����N�*�b��ԋNY^�,�ݜv�z�)��n�{eY�e��N^)��v�˻�����ն�     ��N�   �G�+_)�I�{��C���x��*�M�dQO�7ͤL�u]��M]n��$��L7M���zP�� uS�7�8I֛r���lR�u:MY�eQ��u�u���_w�y��N�����iʬ���Z_$�v��遢I��:I:ESe�2iʲ����kVE�4EYn��z�$���,��N�l���<Iʲ��e�*�f��֧o���*�Ŧ�W�n^M�^���)���_\�yit5/����?���      �
�;    ��Ϸ����k��W�����q�{�WgS��us��ϻEy�t�{WiVU]~���%     ���    ���ߘ�Irg�s      �à��            ��          h	�;           � p          ��           ���          �V�          �
w           ZA�          @+�          h�;           � p          ��           ���          �V�          �
w           ZA�          @+�          h�;           � p          ��           ���          �V�          �
w           ZA�          @+�          h�;           � p          ��           ���          �V�          �
w           ZA�          @+�          h�;           � p          ��           ���          �V�          �
w           ZA�          @+�          h�;           � p          ��           ���          �V�          �
w           ZA�          @+�          h�;           � p          ��           ���          �V�          �
w           ZA�          @+�          h�;           � p          ��           ���          �V�          �
w           ZA�          @+�          h�;           � p          ��           ���          �V�          �
w           ZA�          @+�          h�;           � p          ��           ���          �V�          �
w           ZA�          @+�          h�;           � p          ��           ���          �V�          �
w           ZA�          @+�          h�;           � p          ��           ���          �V�          �
w           ZA�          @+�          h�;           � p          ��           ���          �V�          �
w           ZA�          @+�          h�;           � p          ��           ���          �V�          �
w           ZA�          @+�          h�;           � p          ��           ���          �V�          �
w           ZA�          @+�          h�;           � p          ��           ���          �V�          �
w           ZA�          @+�          h�;           � p          ��           ���          �V�          �
w           ZA�          @+�          h�;           � p          ��           ���          �V�          �
w           ZA�          @+�          h�;           � p          ��           ���          �V�          �
w           ZA�          @+�          h�;           � p          ��           ���          �V�          �
w           ZA�          @+�          h�;           � p          ��           ���          �V�          �
w           ZA�          @+�          h�;           � p          ��           ���          �V�          �
w           ZA�          @+�          h�;           � p          ��           ���   ���k�    ������8      `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap���    IDAT          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          b��,����>�3�6�����m�8�$\�Ans"Ѵ$W)+ը�J�-I����n��3s������q�E���\jc��Հ�D���Rh�-!Q��c�ΜOpS�{�rμ��s��������:��          �N0p          ��          �w           :��          �N0p          ��          �w           :��          �N0p          ��          �w           :��          �N0p          ��          �w           :��          �N0p          ��          �w           :��          �N0p          ��          �w           :��          �N0p          ��          �w           :��          �N0p          ��          �w           :��          �N0p          ��          �w           :��          �N0p          ��          �w           :��          �N0p          ��          �w           :��          �N0p          ��          �w           :��          �N0p          ��          �w           :��          �N0p          ��          �w           :��          �N0p          ��          �w           :��          �N0p          ��          �w           :��      腜� �   ��2p      z!�|^t    �e�      ������;   ��3p      z����    �,w      �/�    �d�      �PJyzt    �e�      �B���   `��      �PJyFt    �e�      �ų�    �,w      �/�Ft     �e�      ��ӎ=��    L��;      �=�Х�    L��;      �����    &��      ��h���    &��      荜�K�    �w      �O^\J��    L��;      �'O��FG    0�      @���G7    0�      @��R�   ���;      �+�    ���      蕜����   ���      �377���    ���;      �;��WE7    0~�      @�l]��;   ��      ����gϞ�FG    0^�      @/UU��    /w      ��~1:    ��2p      �꒥���DG    0>�      @oUU���    ���      ���u��   `Jx�      ������?   �x�      }���     ���      ��u]    `��     ���p�޽�(:   ��3p      z/��/�    �>w      `�d8�4:   ��1p      ��/G    �=�      �T�9���0�   ��3p      ���g��Rt    [g�      L����űc��    l��;      05J)?�����    `k�     ���s>�    ���      ��e���?   ���      Sg4��    ���      ��o7M�S�    l��;      0���    `s�     �i��M��Xt    g�      L���[�    �8w      `j�R������    l��;      0�rUU�::   ��1p      ��/�×FG    pn�      ���9��    ���      ������    ���      3!缸���+�   ��g�      ̊=u��?��    ���      3c4������    |�      ���9?}nn�pt    ߟ�;      0k�YXX�8:   ��2p      f�������    <��;      0sr��xii駣;    �^�     �����(� �,WU��VWWwE�    �(w     �i0�G7 ���ĉ�   ���    8���Zt LBUU����%�    <��    �s�F.�0�J){���W�;    x��;     �TU�� L�+���k�#    0p    `���]p`�UU���p�7�   `��    pN.�0�J)WU���   �Yg�    �9�������+�\�4��;    f��;     ��; 3bw��������C    f��;     �4��	��+N�8qMt   ��2p    ��N�8�`t 씜�[���e�    ���    �s������zt �󪪺euuuWt   ��1p    `�\q`f�R�8y���    ���    ��:  ;���EG    �w     6�w f�yUUݲ���+:   `V�    �Q.�0sJ)W�<y���   �Ya�    �F�0�����FG    �w     6���  r�h4�P]��G�    L;w     6�w f�e���    �v�     lH)�/�  د�m���   �if�    ��TU��� �K)7/--]   0��    ؐ�h��� �Ϩ����   0��    �(���j��@t   �42p    `Cr�.������^   0m�    ؐR�� �󪪺���=�!    ���    ��2p�����{�6�    ���    ��F� �W���4��;    ���;     RU՟G7 @G�wee���    ���    �9}��wRJ�� ��������   �w�     lH]�k��oGw @G�h߾}7EG    ���;     �s��� �R�UMӼ1�   ���    �w xb����tEt   @_�    �� ��ί�������C    ���    ��9���]:77��RJ�   �w     6��b� �m���    �w     6�� 6�MӼ":   �O�    ذ�� �Gv����p8���   ��0p    `�F��� �9O�������O�   �w     6�����REw @��R�(��/�   ��    ذ��Ϥ�\q�M*�\ն���   ��3p    `Sr��  }TJYl���;    ���    �M)��at �T�R�uyy���   ��2p    `S�`[�<�>~����   �"w     6��  ��9s�RJ�   �w     6�E ���m��#    ���    �M)��� �Q�ë�#    ���    �My��H)��; `
���m��dt   @W�    �)u]��93� �����;��yvt   @�    �i���G7 ��(�t�����!    ��    ش���; �����꺞�   �d�    ���F#w �����۷���    �d�    ���� �QJ9ж�Dw    D1p    `�����`BJ)�j����    �    ش#G���ҩ� �R�R�o///�(:   `��    �i9�R��� �b�F��]���ό   �I�     l�ף `�=s0ܵ��rat   �N1p    `Kr��#� f��F������C    v��;     [RJ��� 0J)�ԩS(���   �I3p    `K���jt ̊R�UMӼ5�   `��    ؒ����)�� 0+r�7�m�+�    �d�    ���KJ�Ew �,)���i�+�;    &��    �-+�|5� f� �������!    �`�    ����`�=)�������F�    ���;     �a� 1�VU՝G�}zt   �8�    �e�w��jJ�Dw ��z�3g�]YY�0:   `\�    ز�H)=� 3������p����C    ���    �����  �q�<{���u]�E�    l��;     ���� 0�J)����_)%G�    l��;     ےs6p�nxC�4o��    �w     �emm��RJ��  ���[ڶ�&�   `��    ؖ#G��,�|=� xD)�i���Dw    l��;     ۖs��� ���K)�ٶ�ߋ   �,w     �-���� ��ؕR���m_   ��     l��; tO)eO)宦i�ft   �F�    �msss_I)���  �R�'��y^t   �F�    �mx8��_�; ���9?=�t����s�[    ���    ��(���  <��F�YXX�8:   ���    0.� �a������>u�7�`t   ��1p    `,r�_L)�� �	�����=���O�   �~�    ���Y)���; �s�|4�����g>:   �2p    `l���?� ؐ���w��Ѻ�Ϗ   ���    06��/F7  �������u�;:   �/�    06���� ���j~~��ǎD�    �d�    �]}���3���� `S�?~�#w   ��    ��E  ����Ǐ�\׵?d    ��	     ƪ�r_t �%o������   ��a    ���9��  l�/��ϯ�Rrt   0��    ��>�R�Ft �eol�v%:   �M�     L�}� �����i��#   ��c�    �ؕR�������   `��    0vgϞ�/�4��  �'�|�m��;   ��a�    ��]���N)}%� ؾR�ۚ��.�   ��     LD)�� `l��4Ϳ��    ���;     �s�'� ���m{Ct   0��    ��S�N}.�t2� �R�ی�  �I2p    `"�>�s�tt 0^F�   �$�    0I��  Ư��i�mt   0}�    �����;SJ%� ����   �f�    ��9r�)��Ew  �ֶm-:   ��     Lڝ� ��Rj#w   `\�    ���htWt 0YF�   ���    0Q�\rɗRJ߉�  &�����;   �~3p    `���߿�s�;� ��Rʑ�i�SJ��-   @?�    0q��;� �����˫u]��   6̓     w�ԩ�r�Fw  ;���}��}����   �_�    ����,��� �R�U��󷮮��n   ���    ��s�#� �q�O�<yG]��G�    �`�    ��x��?�RZ��  v�/�ݻ�����'E�    �g�    �����뿝R�|t ��r�?7��^\\��   t��;     ;��rGt �������D�    �e�    ���FI)��  ̏�����   x<�     �#G�|3����  N��o�F�/������   �{�    �Q��ۣ �p/X__�����E�    �b�    ��*�K)�Gw  �~t4ݿ����   �;�    �Q������; �N�d4}fii��!   @7�    ���  �J)WU���pxYt   ��    �WUՇSJg�; �θ(�|_۶/�   b�    �㮹�樂��  :�����ß�   ��    ���  �s.�9rii���!   @w     B���}$��Pt �9TUuw�4':   �y�     �����"���� ���SJ��m��E�    ;��    �0��[� ���]J�m8�):   �9�     �9}��'SJ� t� ��4���   `g�    ��뵔�m� @���b۶��   L��;     �J)��  t_)�H۶��z.�   �w     B:t�k)��Dw  ������ߩ����   `2�    �[� �޸r~~�����}�!   ���    ��rkJ�lt ������xjt   0^�     �;t�П����  z��w���饥���C   ��1p    �J)7G7  �syUU_Z^^�4:   w     :����w���(� ��F_��G�    �g�    @'�u��Rzt �K�?۶�ˢC   ��1p    �3���nJ)�Gw  ���R�=MӼ*:   �:w     :��;�R�7� 譽)���m���   `k�    蔜�M� @��.��6�   l��;     �r��ɏ���8� �A�y�i���!   ���    �)u]���}t �{9��ض�B)%G�    c�    @笯�ߔREw  �WJ9Ҷ�o;vl�   ���;     �s���o�R��  ���?~G]�{�C   �'f�    @'���  L������i��E�    ���    �N���k�N)}=� �*?QJ�������!   ��g�    @'�K)�� �t�9?nn�������   ��    ��htsJ�Dt 0u�z���KKK?   |/w     :�ȑ#'K)�Fw  S��UU}�i�   <��    �N�9�;�T�; ��t^J�Cm����   ��     t����{J�� ���R�۶�Bt   `�    @�R��  L�Rʑ�p�ǎD�   �,3p    ��<�����Gw  �-����Ǐxyy�I�-   0��    輜sI)�zt 0�\__����ʅ�!   0��    �S�N} ��g� ���9���������όn  �Yc�    @/�u�`)e5� �/�7M��   �%�     ��є�C� ��xvJ�KKK/�  �Ya�    @o:t�OSJ�Ew  3�)�����p��!   0�    �R�rJ�Dw  ����'����p���   �v�     �ʡC���s�Tt 0s9�զi��  �if�    @�F��� `&��;۶}_]�s�1   0��    �C�}:���� `6�R��}�>\����   �6�     �R)e)� �]������f8>#�   ���;     �t�������� ̴�9�m��  �ia�    @/�K�y1� �y�)�|�mۗE�   �40p    �����gݖR��� `�=��rO۶��  ��3p    ����߿�t
&    IDATs^��  H)�-�|�m�7G�   @��    �k�v����ҷ�;  RJ�R�o�m��RJ��  �>2p    ��8�p�y%� �/�R�m�����]�-  ��a�޿,;�:��s�+�T�!\�wD��:�E1�E��a �T�9� ��:ҫ��ާ��M@�K&D��`���@�qDְ�QQF���n�Tw�g~ GIwuwU=��z���w��z�Qc�    ��o��,� �u^���z����=J�   �(1p    `�u�݃є�  �O^[[�aii���!   0*�    9�K�+� ����v�}S��{t�   �     ��� C�)���u���!   0��    ^q ��=#�ý^���!   0��    ^q ��I)��z����!   0��    +^q �\J)�m��⪪��  �o�X    `�t�݃9�t ���w���\^U�ɥ[   `��    0�~-"��t �Q�����G���s��!   0,�    ;�n�`D�)� p49��OOO��4��K�   �00p    `,8p`D�u� �xH��u]?�t   �f�    �X��j-"~�t ��+"���zs�C   �$w     ��Ν;+"��t ���R�����K�   @)�     ����������  � E�R�4WU�>   �1    �X�t:�7��  89�]���着��[   `;�    0	�� ����Y333��z���n  ��b�    ���t:WE�5�;  ��J)}���?�t   lw     &�`0X��A� �����`p����K�   �V3p    `"����J)]^� �8��j����zg�  ��d�    ��h�Z����Kw  ��RJ��z��t   lw     &�����"��;  N@J)]�4͛���*   ���    ���n�%"�X� �D�_6;;�����^�   6��;     e~~��)�=�;  NT���333�^t�E��n  ��b�    ��ٱc�%���  ���>��i^:   6��;     g׮]�G��Jw  l���o���I�C   �D�    0�/���Kw  l�S#�C�^o�t   �w     &RJ)�_�t �&99�ty�׫J�   ��2p    `bu�ݛsο]� `��҅u]_ZU�T�   8V�     L�v�}AD,� ��^:;;�������!   p,�    �h�RZ*� ��r�Om��7����n  ��2p    `⥔��\� �-���`pþ}�Y:   6��    �����pk�yw� �-�������z�*   Gc�     ��v����Jw  l�{��>�4�J�   ���    �������  �"�9����z�)   w��     ������d����  [(����u������(   ���     �N��~m���Jw  l����~pee��C   ���    ��YXX�RD��t �6x����MӜQ:   ���;     |���5"n.� ��+�|����cJ�   @��;     |����ʈX/� ���j�����O/   �     p':��E�[Kw  l���`�{�^�e�C   �l�     pZ��k"�Kw  l�����^�W�S�   &��;     ܅���/E��Jw  l��R��i���߿G�   &��;     ���7��  �f/\]]�����=J�   0Y�    ����Z����C�[  ��S���>�w�ޝ�C   ��     p��9_\� ����iyy�{J�   0�    `<xaD|�t @�k�Zk���C   �     �UU}%"^Y� �������~y�   ƛ�;     lP�ӹ2����  �LE����8�J�   0��    �LMM�|D|�t @)9�]MӼ����K�   0~�    ����!"~�t @a?533��������!   �w     8F;w������;  
�������ݻ�t   ���     �����z��ziD��n (�QSSS7�u���!   �w     8�����;  ��}#�M�<�t   ���     �Ӂ^R� `����4�+K�   0��    �8UU��s~ID��n �������*{   ���     N@�۽9�tI� �a�s�u�)�\����V�  ��c�     'huu�5�ץ;  �EJ�9�������{�n  `��    �	���+9�ED.� 0D���v����#J�   0:�    `t��k"�7Jw  ���Z��{����  `4�    �&9|��#�oJw  ��ҽSJ��z��K�   0��    `�\p���s~y� �!tRJ�^�W�  `��    �&�v������  B)�ta]חVU5U:  ��d�     ������E��-� 0�^:33󁥥���!   w     �d\p��F�K""�n ROk��7,--�^:  ��b�     [���\o+� 0��n�oj��K�   0<�    `�LOOϧ�>_� `�= �|}��z�   ���;     l�]�v�/��\� `�����u}N�   �3p    �-���xu��ͥ;  ��tD��i�_(  @Y�     ��#�/JG  ��s�庮߶���c   (��     �X��=�s�وX/� 0~vuu�ʽ{�~K�   ���;     l�n�{c�yo� ��䩩���ݻwg�   ���;     l��V�;  Fģ���n�����C   �>�     �M��:�n�_��n ����5M���!   lw     �F����+� 0BN�9����W�  `��    �6;p���qM� �Ҏ�K�����*[  �1��    �mVU�����/��/�n %9�]333�UUur�   ���;     p�|>����  #�y333׮��ܻt   ���     
Y\\|wD��t �z���ڍM�<�t   ���     
�9�*"��t �zH��u]?�t   ���     
�v�#���V� `�+">����.  ��0p    ��:��E�/��  Q'��.��zU�   N��;     �썈kJw  ���R��i�7WU5U:  ��g�     C�������#⋥[  FU��e333XZZ�-�  ��1p    �!�{�����  qOk��W///߷t   ���     �H��yW����;  F���Z�������!   w     2'�t�|J铥;  F����?����t   g�     Cf׮]������n q���z�/  ���    �ZXX�L��e�;  ��I)����zU�   ���     �T�۽"缿t �H)�뺾�����1   �5w     b</"��t ��x���컪��{�   ;     ���nk�ZsqK� �q�s~���̵�^�>�[   �f�     0�>�s~Y� �1�})����Q:  �;2p    ���v�H)]Z� `�<��n���'�  ���    ��X]]�\� `��W�z���!   |��;     ����nϋ�[J�  ���SJ��z�W�  ��     F�����)��+� 0f�)�_m��⪪l)   
r�    ��Y\\|gJ魥;  �M�y�)��rE�߿[�  �Ie�     #huu�U��  �&����`pu]��V�  `�    �����`0��[  ���眯�����!   ���     F�����9�+� 0�RJ�����~l�  �Ib�     #���^o.� 0��������  ��     0�fgg_7��  S����u]��t  �$0p    �w��j��s�w�[  �T;"��4��9�T:  `��    �����BJ�"b�t ���9��������Q�  `\�    ��X\\�D�yw� �q�R�����+����-�[   Ƒ�;     ��n�{QD��t ��{����MӜQ:  `��    ��i�Z�H)}�t ���Μ�M��ˏ)  0N�    `�,,,ܚs�Ɉ���-  c���V뺺��V:  `\�    ��t:�'"��[  ��lD��i��  �     0�:��UQ��  � �9����zU�  �Qg�     clqq��9�w��  � )�ta]�o��j�t  ��2p    �1�Rʃ��E�[  &ċggg?���4[:  `�    ��۽{�����OF�-�[  &A����v��.���-   ���     &��ݻ�<��3�K�  L��=|���u]{�  �Qb�     ���/"�Jw  L�E�Ǘ���X:  `T�    �9p���r�P� `���j����zg�  �     0A��:t��ץ[  &�I)�߮��եC   ���;     L�׾��_l�Z?��n � ������~UU�   w��     haa�OZ���"b�t ����������N.  0��    `B-,,�AJ��  �'gff�ܻw﷔  6�     0��ҥ�;  &�MMM}�i�3J�   w     �p333��9�t �zT���^����!   ���     &ܹ�{�СCω��*� 0��R�h]�O*  0�    �x�k_�ň�񈸥t ��gD|���͕  (��     ���N��qvD��n �@'��.k�敥C   J2p     ��N�seD���  ��s~C�4�S�  ��    �;�t:{SJo-� 0�rλ��y����w�n  �n�     �7Y]]}UD�X� `�����z����=J�   l'w     ��TUu����Y)�ϗn �`O^[[����?�t  �v1p     ��y�����ώ���[  &أ���KKK�(  ��    ��t���*�|NDJ�  L����O,//?�t  �V3p     ����'".,� 0�Nm��n�晥C   ���;     pT����O)]V� `���s~O��{I�  ��b�     UJ)�ر��q]� �	7�R����_,  ��    �ٵk��V묈���-  .E�/�u��UUM��  �L�     ��-,,|)�����[  ���ξ���߭t  �f1p     �I���l��zfD,� 0�r����ٳ�^�[   6��;     p��gJ��X/� @<nzz�cKKK��  8Q�     �qY\\�@DtKw  �j��7,--=�t  ��0p     �[��ٗRZ)� @DD��n�?�4��  8^�     �	Y]]�O)��t  qj���M�<�t  ��0p     NHUU���OG�M�[  ���Sr����z/)  p��    ����pkD<+">S� ����J)]�����!   ���     ��N�����GĿ�n  ""RJ�¦i.���F  	�     `�����YD�DD�^� ���9��ͪ��K�   ��;     ��:��u9矍�\� ���9?ff�ʕ��{�n  8w     `�u���SJ��  �����~u�׻O�  ��b�     l�����o*� ��K)�ǔҍ�~���[   ;     �efggw��>\� �;x�`0�nyy�1�C   ���;     �e�=��C���gEč�[  ����Z�뗗��Z:  ���     [�����""��t  w0�j��_��sK�   �w     `�u���9?-"�P� �;8)".o����!   �     �6�v��m�ZO��)� ��s�oj�fo�   w     `�,,,|��j���n ��rλ���ժ��I  �b$     ��ZXX�X���X/� ��_5;;������Q�  �L�     ���v��K)��t  �,������߿�KfJ�   ���     (bqqqD�r�  �ԏ�z�W�ٳ�^�C  ��b�     ��t.L)��t  w������[ZZ:�t  09�    ���8��r��.� ����v�}}�4/  Lw     �������� "�+� ��z`����i�C�  `��     �UUu�����"�S�[  �S�圯���)�C  ��f�     �]�vݲ���c��-  ܩ�������[:  _�     ��ؽ{�ߵZ��D�?�n �N���z���  Ɠ�;     0T>ό��[  �S���^�W�  Ə�;     0t:��F�\D*� ��J)�{�^/�J�   ���     J�N�ʈ8;"�K�  p�RJ��iޱ���[  ��`�     �N���ȥ[  �K笮�����߭t  0��    ����tޑs>�t  G���`�+++�(  �6w     `�u�ݕ����  ѓ��֮YYY�w�  `t�     #����Bι_� �#z����uKKK��  F��;     02:�N'����  ѷ������V:  =�     ��H)�3�8�܈���-  љ�V���i��t  0Z�    ��277�~���Dĕ�[  8��r�m��J�   ���     9UU�8p�)��K�  pDߚs�����SK�   ���     IUU}�СC�J)}�t  GtJ�������[:  ~�     �Ⱥ���uǎO�9�Y�  �h:".o��ťC  ��f�     ��]�v��`0xjD|�t  G��9��i���!  ��2p     F��ݻ���j=%"��t  G�r�M�4{K�   ���     �i�ZO��/�n ��rλ�~CUU�+  �8     ��������3"�@�  �ꕧ�r�;���*  w     `�t�ݛs�gE�m�[  8���N9��WVVN*�  w     `�t�ݏD�OD��[  8���s��֮\ZZ�-�  �g�     ��N��8;"�n �~��n_�gϞ{�  �2p     �V��yoJ霈X/� �Q}�����]t�i�C  �r�    ������Μ���� `|��Ç�k���!  @�     ���v�W��^��-  ��s�������  ���;     0��FD.� �ѝ9���z�Y:  �^�     ���t:o����  l�}SJW///?�t  �}�    ����t.N)-��  `C��j����z�_:  ��     ��Y\\���t  �)����yr�  `��     ���V��t  rJD����?�t  ���    ����t^�RZ*� ����>��4�sJ�   [��     �h���KJw  �!�9�w�u���!  ��0p     &ZJ)/..�|D��t  Ҏ�_�����C  ��g�     L����_o)� ���"��u]ϗ  6��;     @|u�s�Η��.+� �����7Msa�  `��     |��������s��.� ��䜫��__�  ��      _����g�y��"⿗n `�^[��%UU��  ���Q     �����w��yN� ��W��̼��+�h�  ���;     ��0r I�|��������(  w     ��077�>;;��K�  �ag8p��UUM�  ���;     ��{�<��煗� FF�������VUur�  ���     �����Ν;�3g?    IDAT�	#w �Q�333����w+  l��;     �� ������_y�%�̔  6��     `��� FOJ�o���_ZZ�-�  ��;     �10r =9�'NMM]���r��-  ���     ##w �ѓs~����5�~���-  �]3p     8F�  #�9����s��!  ��3p     8N�6rO)]V� ���9����G����-  �73p     8sss�g�q��� ���䜯۷o��J�   wd�     p��� FOJ�����,--ݿt  ���     6��; �H��v�}M��@�  ��     6��������#❥[  ذG�k���N/  �     l����ܹ�#��[  ذ����������!  0��     6��������"��J�  �ag�k���R:  &��;     �H)����WEį�n `cr�;[�ֵ���+�  ���     `�|m����E�[  ذ3Z����~�Q�C  `�     l�����#b�t  v�`0�H]��Q:  &��;     �6�t:�s���  `���z�  ���;     �6�v�KF�  #�>���#w  �>�      ۨ��.ED�t  v��`pu]��Q:  &��;     �6�t:MD���ȥ[  ؐ�"�#w  �z�      t:�7�ύ�A�  6䴈�f߾}�,  ���     ��n�{i����8\� �9m}}��  ���;     @A�n�2#w ��r��������� �qd�     PX�۽<����8T� �9}0\������!  0n�     �������ϊ��J�  �!��Z-#w  �d�      C���~0���0r g���kz�ރJ�  ��0p     "�n���V���Z� ���9�L)}l߾}.�  ���     `�,,,|,"�_*� ���1�5r �g�     0�:����~$��O�[  8�����`pm��{P�  e�      Cjqq�SJO���-� ���w�Z��� ��3p     b�N����'D�_�n ��r�;SJ��۷[  `�     ����ϵ��'Fğ�n `C�\__���;  ;w     �0??�����'G��*� ������~U��@�  %�      #�����v���qc�  6䡃���}��ݯt  �
w     �2??���S"���-  l�����?�gϞ{� �Q`�     0b�������K)��t  �]�������� �ag�     0�v��u����\D��t  ��`�������!  0��     FTUUk;w�<;"�V� �y���ԕ�\r�L�  V�      #lnnn}qq�%)���-  ]����z�{��:�t  #w ���w�_�_u�ǿ��Nwb�AV�b���(0K��@�$�X���t��:���tg	��hb�9�:�D	a!� � 
3(K�AD.	*	]!����y D I�/U�������>ko    �\J)w:��9�~�  �Y333o��꫷� �Qc�     0RJ���:缫t  ��܃��i�-�C  `��     L����RJ݈ȥ[  8���SN<���4Mc�  ��8     �0�nw9"���[  8���E333�6r �op     L���^�s~zD|�t  ��9���W��  �Q`�     0���������t  ��s�x0�-�  ��     L�n���#�̈�b�  -缳��_V�  J2p     �pUU�ED��\� �{��~�i�  (��     `
TU���v�1�[  �G������  P��;     ��XXX��p8<5"�_�  -��4~�t  l6w     �)�����V�������-  R�9�|0<�t  l&w     �)��t��s>3����-  R+�|�`0���!  �Y�     �P]׷�߿�	qc�  ��s~�����K�  �f0p     �RM����{fJ�ե[  8��9�7���ǔ ��f�     0�����:���s���-  ܽ���D��������-  ���     �\J)�u]�w�n ����j��x0�H�  �(�      DDD]�K)�Eİt  w�~9�w,--�T:  6��;      w�v���s���8X� ����v����/��>�C  `��     �꺾>��Ԉ��t  w�Ƕn���k��f�t  �'w      ���-������t  w둷�v��7Ms|�  X/�      ܥ�����j��T� ��u�������R:  փ�;      w����]��>5"��t  w�333�5Mc ��s�     pH�޲e�i)��n �n�����U�#  �X�     p�v�����?����;K�  p�r�������  �ca�     �aپ}������7�n �n]6:�#  �h�     pؚ�9077wa����-  ܵ�s0�b�  8�      �������_�s�U� ���rίO+  G��     ��R��R���1,� ���s���ٳ��!  p$�     8ju]�<"�K�  p'[[������C  �p�     pL���ݔ�y��t  w����������!  p8�     8f�n�Eę���-  |���}[��;����(�  ���     �uQU�_����"�3�[  ��>x��ۮ�暙�!  p(�      ���������>&">V� ��R���n��-M�l-�  w��     �u�k׮�[��)���-  �ə333��S�  �+�      ��N������-  ���-//�z�  �+�      l���o]YYybD\W� ��s����v��  ��f�     ��i�f���>/�|Y�  �SJi0~�t  |;w      6TJ)�u�D�Έ� �ߵrί���g� �o1p     `STUuUD<+"�n �[#��={�<�t  D�     �����ݜ�y���-  ��{[�������K�  ��;      �����D���-  �ᤵ��w�z��� `��     �骪�`��Q���-  ���)�?��z'� `z�     PD]ןڲe˩)��n �?�Rzc�4[J�  0��     (f�Ν�?���O�9�Q�  �p��'����s* ��1p     ���۷��z�O��7�n �RJ����Jw  0}�     (�i�+++���,� �7��^���_X� ��b�     �Hh�f��v"bgDK�  /O, ��0p     `�TUuUJ��q�t  ��9�~Ϟ=/ �t0p     `�t����Ϗ���[  ��V����`���!  L>w      FR]��n�Zg���t  qR����\s�L�  &��;      #���|`˖-�����n  ~�m��k�fK�  &��;      #maa�89"�_� �8ovv��JG  0��     y�^z�-9�#��[  �]����~�t  ���     ��P���sssOJ)��t  ����O- ��1p     `l��ϯu:��/+� 0�Z���`��!  Lw      �JJ)�uݤ����{  ��	���{�����!  Lw      �R�۽.������J�  L���}SJp�W|_�  &��;      c���u8��s���-  �*���[�lys�4[K�  0��     ku]�y������-  �*�t����+Jw  0��     {��������>T� `��B�߿�t  ���     ��������?��xG� �)�k����  �/w      &����WVVV��Rzu� �)�rί�+ �x2p     `�4M���t��s��t ��ښs�a0�H�  Ə�;      '���n"bGD�  L���ߺw��{� `��     0����͈xZD�V� `
=tmmm_�4[J�  0>�     �hUU�e8�_*� 0�Ξ��핎  `|�     0����j=2">^� `��w���_*� �x0p     `*t:������t �z�����#  }�      L�����E�c#�m�S  ��q���M{��}P�  F��;      S���[��果s���-  S�>kkk����N, ��2p     `���ϯ�u������=  S�a�V�uM��- p��      L����J)=3"�^� `Z䜟233��  �&w      �Z�۽!�|AD|�t �yI��{f�  F��;      S�����Z�G��n.� 0%RJ�~��S�C  -�      �N��VWWO���*� 0%N���,--�T: ��a�      �t�%���	'�pZD��t ��8��n�x��Wo+ �h0p     �o�}������'��^U� `J�|���t  ���      �K�4��N�9��J�  L��ҳ�A�t  ��     �]H)庮���/F���=  �.����t  e�     �!�u���� "�Z� `µr��///�X�  �1p     �{PUջ"⌈�\� �	7;�|�W|_�  �0p     ��PU�����9珔n �p9����۷�]: ��g�      �iaa�ӫ����9��t ��;��o~i�  6��;      �ݻwy۶m�F�J�  L���z����  `s�     �ڱc���n��rΗ�n �`)�t����K�  �y�     �(��r]�MD<?"V�  L�{�����z'� `s�     �1���期�R�Z� �	��)�W��  `s�     �1����SJ���/�n �P�����  `��     �:�t:h��'G�?�n �P�={��Z: ��e�      �daa�8%"�W� `�j��---�T: ��c�      ���K/�eee���W� `ݿ�n��4���!  lw      XgM�|}nn�gSJ//� 0�N���]* ��0p     �0??���v_;#bX� `��w�g��  `��     ���ꪔ�|D|�t �$�9�b0<�t  ���      6X��}S�����b� �	rB���{��w�  ֏�;      l�����n�O���J�  L������N�4vP  �a      �daa�#�v�����-  �	����KG  �>�     `-,,|6�|jD��t ���9�j��?�t  ���      6Y]׷���<%�|m� �	ъ������ ���     @MӬ�u����=  �>qC�4[K�  p��     �����J)�G�m�[  &�O���.��  ���     @a�n�M9�3s��Z� `���{��j�  ���;      ����ߟs>9"��t ��K��{�>�t  G��      F����'8pJD��t �����������m�C  82�      0B.���[VVVΎ�7�n g)��<p�@�t  G��      FL�4_�v��/+� 0�^���~�t  ���      FPJ)�u�D�ΈX+� 0�RJ�XZZzh�  ��;      ������9�LJ�k�[  ��l��~C�4Ǘ ���     ������)��E��K�  ��G����) �=3p     �1��t>�s>9">Z� `L]����\: �C3p     �1Q���<xJ����[  �P������K�  p��     `��޽��۶m;7�t}� �1�})���۷�]: ��f�      cfǎ�w:��rΗ�n 79�S?���J�  ;      ���R��I)=7"�� '9��z�3Jw  pg�      0ƺ��uqAD|�t �i��~����  ���;      ������j��)� 0F~0��ڜs* ��3p     �	��t>���������-  �"�t�`0��t  ���      &Į]�n^[[;%"�Q� `�����JG  ��      0A.���+++O��W�n �r��///�P:  w      �8MӬVU����ȥ{  ���W��  ��      &V]�K�q�t �����.( 0��     `�UU�ڜ�y�o�[  F\J)]w�W�@� �if�      �����Z��D�M�[  F��VWW_�sN�C  ���;      L�N��w�v���`� �w����/��  �V�      0%>�s>="�V� `�-����T: `�     ����ֹ��'G�o�n U9��I)�n�4[K�  Lw      �2���kUUm���1,� 0�r��uvv�)� 0m�     `JUUuUJi>"n+� 0�rΗ����Jw  Lw      �b�n�M���܈��t �jEī{�މ�C  ���;      L����?������n A��^� �ia�      ����'Z��)�'�[  FMJ酃����  ���      ���N��[���R��t ��I9�W-//���!  ���      �Î;n�t:�/+� 0bN��* 0��     ��R�u]7)��F���=  #䩽^#  &��;      p����u9��#�+�[  FEJ���Jw  L*w      �n�u��V�ujD|�t ����p8|E� �Ie�      R���p��~d��/K�  ��������9�;  &��;      p�>����N 	9�+��Jw  Lw      ��u}����S#�7K�  ��{��W��  �4�      �a���_��jGD쌈��=  %�������.� 0I�     �#VU�U�����J�  v������  ��      �Q���-qJD�S� ����n�_Q: `R�      G����M��zTD�u� ��.����. 0	�     �c��t���n?.����-  ]����C�#  Ɲ�;      p��m۶m�F��[  
�W�����  ���      X;v츽��>#"z�[  
y�`0xF� �qf�      ���R��j1"vFİt �f�9��ꫯ�o� �qe�      �������gD��K�  l��?p��m  ���;      �!���1�|AD|�t �&{��={�) 0��     �S��{Z�֩�O�[  6S��z�5�\3S� `��      ���|��n�-� �����}��  ���      �p�n�Z�����n �,)���^���  ���      ��N�K[�n=+"n,� �IZ)�k�����J�  �w      `��ر�����gF�+K�  l�_YYY, 0.�     �M5??�VU�rλ""�� �h9�,--=�t �80p      ���z)"~!"�n �`۶l�ru� �q`�      SU�k#₈�_� `#����z�,� 0��     ����zWD�_(� ��RJ{���{��  ���      (����h��'G��K�  l������Z� �Qf�      �����Onٲ�Ԉ�`� ������?]: `T�      #c�Ν��9��Rzg� ����j�fK� �Qd�      ����oݿ�"��-  �'N<�ċKG  �"w      `�4Ms`nn�ҫK�  l��ү.--�P� �Qc�      ������N�����e�[  6�l����  5�      ��J)庮����p �z����疎  �ޤ  �IDAT%�      �ȫ�ꪈxvD��n XO9��^{�q�;  F��;      0��z]J�iq[� ���R������(� 0*�     ����v��j�΋���n XG/[^^���  ���      +�N�qFD|�t �:��K�#  F��;      0v���`��>9">Q� `��\��{l� ���     �������v�}jD|�t �zH)���k�=�t @I�      ��ZXX����O����n X?�����  (��      k�w���	'�pND��t �:����ݯt @)�      ��۾}�������t �1�WD�j� �R�     ���4́�����9_[� �X������~�t @	�      �Ę��_����9�]�[  �A;�te� ��     ��S��RD숈a� ����~����  ���      �HUU�fJ��q�t �Q\}���JG  l&w      `bu��ק����n 8
:x���KG  l&w      `�u�ݷ��K�  ���K���s��  ���      �xu]���8?"�R8 �Hͦ���  ���      �
UU���j���n 8)���z��(� ��     ����t���n��R� ��SJ{JG  lw      `�,,,|$�����T� �#pn��?�t �F3p      �N]ןZ]]}lD|�t ��5Mc� L4�      0�v��u�p8<-">\� �0=lvv���  ��      �Z����;x�����-  �#�|y�4�S� `��      Sm���_^]]='"�o� ����333��  �(�      ��۵k�Wr��DĻJ�  �ݗ_~�}JG  lw      �����֭[�>!"�R� ��{۶m�R: `#�      |ӎ;n_YYyFD�P� �Pr�/Z^^~p� ��f�      �m��9077wa��wJ�  �֜�e�#  ֛�;      �w���_���9qU� ���s~�`0xX� ��d�      pRJ����9��Q� �n�"�+� �D1p      8���_�s�U� �䜟���N.� �^�      �A]�K)��#"�n �n)��(�  �^�      C�۽&"^��-  ���`pf� ��`�      p���ze���#b�t ���9_�sN�;  ���;      �������0"�n �6?����X: �X�      ���nL)=9"�^� �[RJ��4�M 0�3       G����aJ�ia� ���233sa� �ca�      p������'E�m�[  ��eM�l) p��      �����;#���R�  "233��  G��      �UU�'q^D�/� /۷o_�t ��0p      XUU�o8�_-� L���t�M^q ƒ�;      �:Y\\���8#"�T� �n)��+� �82p      XGUU}p8���n ��Cn�����  G��      `�-..~h8�_,� L���K��� Ɗ�      `,..�u��>-">W� �N)�=���� �w      ���������- ��z�W��q�p      �@u]�m���0r 
��+�O/� p��      6X]��G�gK�  �'�ti�9��  8�       �����F�a� l���sJG  w      �Mb� ��s�]� �p�      l"#w �����{��yt� �{b�      �ɪ��������� �D�VkW� �{b�      P�%�\�1#w `�]0Q: �P�      
1r 6Y���t ���      d� l���3���\� ���      v�%�|,"Ί�ϗn &^{mm�+� ��2p      UU��������- �dK)=��+����  w��      `D\r�%k�Z�D�K�  m����KG  �w      ���t>�R:+"n)� L��p�}yy���  ���      `�t�ݿ�gEėJ�  �)�tߵ���Jw  |7w      �����������r� `2���M�ؐ #�q      0�?�s� "��n &�Cggg_: ���      �����?ϋ���- ���9wK7  |;w      �����ga� l�3��#JG  |��;      ����}9�D�m�[ ��2;�  ���      `L�u��V��Ԉ��t 09RJ�XZZ:�t @��;      �X�t:�j��F� ��9��j�R� �w      ����t�(�|aD��n &CJ�M�l-� `�      0��~sD\k�[ ��p�������  0p      SUU�ύ�a� `"\\:  ��      `�UU�ڔҎ� �D8eyy�'KG  ���      `�u��kr��; ��7�t 0��      &@]�W�/+� ��/������  ���;      ���뺉��(� ���n���� ��2p      � UU��9/��  �ڋ����. L'w      �	SUU�)� ���t�M�/ L'w      �	�R�+++�K)]_� O�V��� ��d�      0���>�xVD��v���һ����=g;���"b
�DEH�1@�L�<�"�5�m�Rim7D2t�9�L��i4���.	A�J�bB�4���D"B�B[���ݝ=��B��>��u�s^�������'�_f�  ӧ���[n���� ��1p      �Q{��/,,\�n �Ύ�d�� `��      ̰���c�^owD|2� �.��ko��~v 0_�      f�`0x`aa�qgv 0=j���}��gw  ���      `,//�����%��/g�  ӣ��]��  �w      �9������d�҈�;� ��:t�й� ��0p      �#�����z��Dķ�[ ����ĉ�ώ  懁;      ��_-��zD|7� �R���ZKv 0�      ��p8�b����X�n :�<��� `>�      ̩�i>Sk�,"�n ������ `>�      ̱�in��^'�[ ���m۝� ��3p      �sM��u)�1�n :k���⫲# ��g�      @���R��; ����zWe7  ���      ����﮵�-� �Z�8��� `��      �CMӴ��� ��z�~��� �l3p      �!����� @']�  �6w       �m����ҕ��� �s�s�-�<?; �]�       <�޽{7���k"�� �[j��� [��      �G������Z��� t�d2��m�� �l2p      �Q�F���L&/-�|=� �R�S�9�_��  f��;       �iuu��Z�%qv �Wd  ���      ��5�����]��- @'��#G�� �w       N�`0�l�uwD�n ������˲# ��c�      �Ik���k�o��Iv ����  `��      pJ�����:��  r�Z_ٶ��� `��      pʚ�9���  R������ �l1p      ���Ո���  O�׻"� �-�       ��RJ]__�.">�� 䨵^r�ȑ]� ��0p      വm{|<�g�  )�>v�إ� ��0p      ����������G���- ��+���n  f��;       gl߾}���z/��~'� �v��m{vv 0�      �����~�7"�hv ���YZZzqv 0�      �4��೥�+"�Dv �}j��� ��`�      ��������  ��em��Ȏ  ���;       �n4������ ��y�����# ��g�      ���Fo���gw  ۣ����n  ���;       [��R����F�ǳ[ ��Wk�]k-� �t3p      `��ݻwc<�&"��� l��:��� `��      ��VWW������ `kM&�K� ��f�      ��[]]��Z���� `K� g��      �m�4͗z��q"� �2/8|��OeG  ���      �m3>o��  �Lo<�,; �^�       l��h���xGv �5j��d7  ���      �m7WK)�fw  [�em��Ȏ  ���;       ۮ�R��֮��Og�  ���;w���� `:�      ��m��?�ʈ��� `s���K� ��d�      @�����7�L.��~'� �<�֗g7  ���      �T+++_+��:"�e�  ��xFv 0}�      H7�>Yk�:"jv �9����� ��1p      �������� ��1p N��;       �1����  6ŋk�%; �.�       tF)��z�k"�3�- �;�����Ύ  ���;       �2�L&���od�  g���  `��      �9+++ߚL&�����- ��+�� ���      �NZYY�B��ʈ�d�  ����km����  ���;       ��4�Gj���� �������gG  ���      �Nk��"�}� �i�8;  ��       t���J)���  N]��� 8i�       t����cǎ]_�n N�/�m�� Lw       �������������g�  �䉋���ˎ  ���;       Sc߾}_.��6"��- ��+��(� ��       L��p�7�?� 8%/�  ���;       Sg4�q)��� ऽ�m[{5 �q9       �Jkkk�D�� �Iy�]��� t��;       S�m�O�8���vv ��&�ɋ� ��3p      `j�p�_/�쎈��- �c+�� ���      ��6?]J�>� xl��_�n  ���      ��7����  �3n����# �n3p      `&,--����� �����bv �m�       ̄�{�n�u�Y�G�7�[ �G���  ���      ��_��R.+�� � xD� �c2p      `�����Z���  ����n���� t��;       3g4}0"fw  s�=����� ���      �I��jD�]v �0/�  ���      ���gϞq���"��� �!��Ge�      ��j��۵�WGı� ����Ge�      �Lk��3��av �J)�m{vv �M�       ̼�p��Z��; ���8kqq�� ���      ��~��R��; ��R�/d7  �d�      �\�R.���e� ����>7� �&w       ��`0�j)�ʈ�d� �<+�\��  t��;       se8~4"ޞ� s��k�%; �w       �����[j��� �9�t���gfG  �c�      ��i�v���_we� ��:q��E� @��      0����qyD�n�y������  t��;       sk4�Qkew ���� xw       �Z�4ew ����� c�      ����{#�+� 0g�y�ȑ]� @��      0�VWW�z���"�Xv ̑����� �[�       "��?�ZW�; `��Z���  t��;       ���i�Dć�; `^�R���0p      ���������; `�� �8w       �����^D\ǳ[ `� a�       ?f4�Qk]�� �9�3m��Ȏ  ���       �h4zg)�#� 0�v��uav ��       �J)���]we� �,����n  ���       ž}���G��� �U����n  ���       �h4�#"ޒ� 3�� �!w       x���7G��� 0�~6;  �w       xm�Nz���#�� �5��� ��0p      ��0���zmv ̚Z��۶]��  ���       NR�4)��Iv ̘�Ν;�ˎ  ���       N�d2ysD�[v ̒~�av ��       p
��9�����- 0+j���n  ���       N�h4����fw ����^��  t��;       ���G���۳; `�R.�n  ���       NC۶��x|UDܟ� 3��� @7�      �iZ]]�7"��� �pav  ��       pF�ч#��� 0��m����  ��;       ���x�戸+� �Xyғ����  ��;       ����յ�dreDL�[ `Zmll���  �3p      �M����Rʻ�; `Z�z=w ��       6���ڍ�� �R� ��;       l��mPk��g� ��)�� �       �����ǈ8�� Ӧ����  ��;       l����ߏ��� �i�; a�       �nyy�X)媈��n�iQk5p �      `+����Zߞ� S�� 0p      ��r��ћ"��� �O9r���# �\�       �Eڶ=Qk�:"�g� �(<��S�# �\�       ������R�M� 0z��Of7  ��      `����(�|.� ���; �9w       �bm۞���#b#� ����=%� �e�       �`8~����� ��d�; �9w       �&G�}kD|-� :�� 朁;       l��mPk�."jv tQ)�� 朁;       l��in��~0� :�� 朁;       l�����#��� �A� 0��      `��߿���ew @���3p      �����K)�� c� s��       ��Z����� 营�   ��;       $�F��Rޖ� ��  �2p      �D�wޡ��3� :�� 朁;       $ڳg�8"��� �'�ZKv ���       ��F�;"�O�; �z�:;; �c�       p���"�� �6�L� �<�       ���￯��fw @��3p      ������_�� �d� 0��      �#���3�L&o���� ��`��      @����|����� �Rk5p�9f�       �cǎ��X�� ��^ogv ���       :f߾}�,�ܔ� Ivd  y�      �����Gė�; `�M&�~v ���       :�m����; `��z=�`��      @G��O�Z�*� �S��� 昁;       t[ǲ# `��R�� @w       谦i�*��'� ��� 0��      ��?~SDܟ� ۡ�j� s��       :��o�nD�#� �C)���  �1p      �)���~����� �>��3p      �)ж탓ɤ�� ��Vk5p�9��<�P����    IEND�B`�PK
      RZ���͗  �  /   images/cc0ca695-66e1-46bc-a2f3-28706ce884b5.png�PNG

   IHDR   d   �   ��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  $IDATx��	�U��������sgr'$�!�Ka��
쪫�9d�#"GP!�7�D�]%A���]9Vv]EvA��H"1w&�$s�Y�u���Wݓ���g�z�z��_^���z���}ǻ�T����
�eR�2�q�T��L�@\&U .�*�I�ˤ
�eR�2�q�T��L�@\&U .�*�I�ˤ
�eR�2�q�T��L�@\&U .�*�I�ˤ
�eR�2�q����nOA"�@��:���8�wz�؉���c:�0���ւ�B�˸���j�i �` ф]�	`b���cZD2��6_�� 
@�'VC � �;8|�F����>���<@c
�w$�;Ρ[u2R jE@X� k��r2B��0���@������K�Ѕr!�B@o��;�4���v:z8|�<�ˇ��C�Ș ��6M�A-�,j��܄��yX��G�8��)פ��$
NG���Ŵ�,ؠz�.�����fO����l5�A��&��)+�ϯKB4ʥ)�D��s��O`+��JE���-�T	�Lt��؎�3LOc�Qj�1*������ȧoҠ��6��ԈE����@�c�d�Sb坓�h%�u.�՘�#���14{pŗHc�xC �&����$��O��VD�J��X�뀜2���O��#0��\�l��.L��c6%��A�N3X�A�O�u��8
�ʛ5�����!��������Ř0�*�$��#�SIaii�!�'+�cd�|�r������1�I�(2�R����|�q�(��dK�(ɋm�kX׀m>ӈ���(�Ƀ^/c�;�q��2�z"�H�p�EϾ~ �˹��')�>ڍ�r
Z?�&� ��0����f��އ__�F(�x���(��/d�ܙ��`��Y�]�D��K�?*S#i�wٮ=p��y�	�zM
���_)���������n�A+
�H�wc~�a�,��Ib��s����;pXdv�ci�Qa*}M�0�?�i�\��Zr3�>��	��P�ϯ���Tưa�Ş��n~=��a�:�	�J�,ut�`��r�5}&S�`�͜�x��eio��JS ��-���Q��˧Q��+���ʨ�\y�&��}�K�0�w�.<�*���-�;����l7�4<R*�}4.�4MS����u"O�� [~
N��<�l��=1ab���LP>��������	�MF�����#얎�5S��`�V���V����a^2����۬�� l�⹗���iL]�����)9M!Ɂ��@��n%����dk���r	jGY���ף��
HO�}�Ma�|l���LQE��2��<�T�Tl�ԂŢy�K�E���bF,9({�́VS_0�{O;�Зpl����³�����_�7�j�^,��~�m�ǺW?b ��I������h���ʟ���w�TB� (�y�r�՞��bhn��:��A�ݹ�Jm�9�y���y��9#�rޙJ�1v��7��s܊���k^�/��M��=vPF�uIh��S��D3ƅ�(ali,�RH���\��\	&����-�D($�
����[���+�М��k4:��3�P&c��G��/�@^<�;x}��kw�Ѯ��2" �Q���j�=p��>�M>��i��9�B!'�?�,|�E3�i 
��
4t���Lp���'��"<:�w���~�[3���˛�\�`�oE kф�U��x��hI�@���,tw�C�j��C��*j}~t�X��LjF���Gx��ؒ_x�L�/p"&�N*Er/��L
on`*:l�����Ңh�̓��
��s4��1�����^J�]�(���)��:ہw�\=Ԅc��j����^�}��A�#�tZNb��)�Ǿ�`���ܒH��5�Ӓ���x�]Q{�=���}�+��ؼ��[j�d���Nێ���֝3Y}�!�Fm��i�H�LV����C�a�szY��KQ@:z�/n��K���A��JQM�*	���63��Ud��r5�_~� b�A!�>͵�~���/����o�WK��jK��>���w������#����@B0�|��� ��+����z�t�����2,��nKA2)�<�	��ى�AY��}����Z*i����z$t=AԒ�������ۭa��4fځ\�0N�+H��7��R�x(�'xd�*@3���hV�w���_K�}�
�-�a��2��)Ǫ/���@���[f1�5�v��QW���_���t��؝Tʚٰ@(�B(4fEb��� P�<f|� 	��hL�o`4E*K��y���͋���rɐ@���.-j��\�8
�PIgNc���!fBع[h�)�0�ȉ����Qh�d9eH =�ޱ�e��G':�T�^�\�p�<�`�ˀ`�k�t'ƫ�I�lͯ	ɩߎrf4$�Y� ���� }+;K�0
2.���
���ҥvT.2��x���r��8lGF�����aC�'z��ȊJ�Ԃ׽�skS���.�b�!����⫌�f�T;����P��̕���P�L���M�K�������Q˨� $47��	HJ���J��:���S��C�Z��ђ� hկ�3t5�8�/���8H$;G_6�5@�86l�d�wC6
�t�k��ޔK��ul�?c��
�+P��2^�k�VŖ*�I�ˤ
�e2�0���d!�k"�ID��z���F
Uů3�1 4vRn ��/��y�C+��W#hɉ�<ɤ����}��v�q��!A�`���@�L2���l�S�;��_��^_]<��7��E82�=�cN1��ߍ}ղ !;m5���ZT�L�^<�t�x#Z 45�w�� ��IA�g���v
W��@�Okq:�)\0{Y`.�_$OM��v�q�&�9l2_�xk]Zk�a.�t�e<��]S�����?P�`&�0PLQ#�V�J�p'瀠��h1��:��`(�� �P���	F*y�&�8\.�tTC�mH�`(�&2��BZ�=���*@&@?C[t�h����`�FZ�&b��Bf *�3��{��	�ad�=�D�`3z72S�@��s���b�[C������f!LVIsc
�6?����>_}�=�E�!�C�MTV(�PxV�?����a�<����`�����g%=���a�!�B%�8c�ah<ֳ��43*�@$��[_pz���Y�呝�=���dl_�ihJn��r��������{`
�%�Æ��h$�Ƨ���4��T�%4�o�T|O���j�� q=	�ט	�Z
n�!�dA2�/�g��� ��1 �p��0z��I�F�ߧ��Fׄ�A��쌠c�C�D�@x 
�;�Jf�^'`�P�D� B���:5Mk����q���a2�q�#�!o`@;�Y�3�!i������o�� ����i9�h=h�����Љ�S����Q��fJX�y��έva�=�A�`�z�������NKI�0TL�䂁��`��i�Hsf$��86X�=��"Zی����(���l�*��y���ܴxP�V�
~NkivqO�_��Og\zm�����~GĲ��$l���[��T<ܠ�ܢ����8_��a��Ք����+����p&��{�O)��`b4@H�}��:��Qs9GV��Q��^�_����(V��:R��k��Ydt����h�v�t�M[�v��nY<@���W�L��WЧ|c�Vݘ������F
�Q!ar��6>�b�{��Q�������wy�t$@��2����1�6�%d��L�I�=^�W��[я^8�ǭh �
�FN�K�(�j�eU�O�}�|&O?Xz�U<��^��2O|��;����TԒ�#���3C�������ߘ²�a �ȳ�����+upB���I!���7H;ʸ!��BZ���������/��DF���P�&e.o(��2e�8���7�/[���Pڳ��q�|�uřkFC�S� >�X�u����٩S'۲`�6ی���+6V2�osC�~dX ��ľ���+��3@^�=�b���=��s>�1�a�E�{%mh� �� ��g�ް���K�YUXvK�[��KO�yq{y)�,5h��s�cT�Bˁ���L�l?Eo4�4dN)��<s�^�<a�pj��r�p����A�jO�Y�D��ePM���b�<�MF򖞎���O�!,k�8/3�L@7�xhk^��v��4�6y�{�y ��Z�¤&�֛L��&�(�a̙��ç`w(c05 b↾�]�aʵ|��+|�����E��Ĝ�Z�Z��0z+�[;`�4$�2*��#4�ȝ�A��9�S�@�*?�qb���cT�>^:���G�\ZB�Ђ�~�C�m�� Y!�Ԙ?c�wH�whi�Й�����x����K���I�����'�Lx�E՛H� �����;�{�ӫ3�:),�춳@c=XG�gfd\*�T� ���;���ǾN��u�fyG,#B��]���i'���7c��FE���G&z0Y�A*с�_�O��ה���|H0�p./��W����ff���L����'Yp���"��/'5�Vr�u3�+��Hf]�|ޔ�Ӄ#9g~��'F'>��� � Z��������!�P��5M{�h;�˯	q�vč&��4�����d�J��@���3�L�U�AUO��.8�**��-�^�@���='#�x���ϥ{�1�
�J�X�Ld�85�~??�講V�?�řյE��N��'���# ���gqV_k��C>/���h�\���i(�x_
a�����f��_���~ҎH�9�0°W�����C �<g��Ogl���$�B�����"7G:�lF�}n[��<h_������xw�ACY>l�ku�u��~f�s{DF����!��M�� ��%!�I<g�¤�Ph�����P[�!"��Kp�0ڡ�@D}+n��1K���6dk��'�~��)���*��sBfz�@ڰ��H�rdR*_F�ފZ=����͚���B�D�zT��1X��1
���cĢ�F�rޙ���f@G���';���cZ�B�N�p�Bkb��@�ZBdM-E��4)0c����}�F�����wP�ώ� p���ա�����:����rT}f��HZ�|Mmb��] ��) ���+�҅�-D3ڭsj�����v���4�;j��tQ���}e�Jn�� �I����847�P_���e���t1sg18xX������1�N�t!��0�젣�꜏a���ЉǓ���+�Ewf�;SEPH[�<$���xg��Wb�[d�뙬�`�aRa�tt]@"iA4nAO̒ﵴ�g�2j���b��D�
�P�~�^����sٱ�+�d9��e�y?�4�]�q��	8���
�	�Y�@?O����%�6��0���G���p++���yi�:Q`�U҅�6�����^0�]{-x}'�ۻ�R-3̜����I�>�W��:[�,9U, a3 g+t,:7���9��1�����+^z��I����6e��[Hm8xD�f��+
�FŬ�S�$������s��ď��)m���>t�A?�^�uô:�1�;�%���`V�
��%^|Ղ]{;��`ˤy��:�&iꠡ����(v%�|�!�7UZ�Ya���u*l��N��P��$a��GH(^�8�v#��������^{
<��|;���!��bC	 �%��a�|���C�B�:^�1�C�%��dZr�ۻ��:v`��.��hj�W��G���K�#MJ�tJd�2h�R����h\�'���5������HF0�g��^B�B{�tKO?������`��I������Ν>�=����.2�dsB�)2�����Q���ĮhnK:�&bok�'�n�A�Z<�0��X.�r9z����5#��{�~-C��#����o�,:�%�uÝiX2���Vk�u�w���4�
�uؒG4�ܻR9q��\���J�`����$4&z?�8=����~��p��,�����#��w�znN��K<p�=F5�YO65�o����<�0�il�gSr�u�Vx=bFQ	
f2�e�Ӱ�2?":OF�1|�{d��w��x�I�k�"�?l7�)b�c�W���y�+`��0��������I3�V�c\�Q�Z�c�,��A(:,]ğ��"��ǟ2.@Ǽ]��B�~��⎝pd܄���
�Z���~dLΉwEU�ڨ;:65R)i��#����oM�b ش9C��/������ ���5�!�5���ؓ��p>��
�������w>���sW5�d���iMt�(���$��OÖ"����ûzM���᰺�H��V8w�kKN�㱹�kA8���>YQr�r}��!��W" ܞ�a&F[	��As�>h��A_�\�����w��K/O��:<���^�h��͜[6aÆ o�Ô�&%�B�P>�T�2���BOr�N�d��0P��&+V���-�d�����%���jBm�����&�fZ
6�6���֬YO�{dv�2Yi � 7�놐�fԿ%��?��h*�����e�w'�ǰuO���~����	�c�3���,��!|�[����8��Q�{b$��� lM��ʸ/�ow�V����GMA���̖�x���������V��3�sH�o�n�7������	��pJ�s�x��k��.����d�7�J�q��k�i�
-ULk�/���E��@���&��W��]���4�i=��=��Y��@Bx�x`���&���d�*�I�ˤ
�eR�2�q�T��L�@\&U .�*�I�ˤ
�eR�2�q�T��L�@\&��kW�MV Ksoh��<q�LV ��/0�}p�J���	���c�+�|n�R�@���S1=����f7@�t oc���0��Y<��j�]�?�P*H���..�W!��� ����R�@H�Ҁ�|
S�O�8��� �IL/c:����_a�;L���R�@��6ث�^k1�ځ���1}�k��XC�X �,��a��皇�7����}1�P*H���|�JL�;pj�'�m䳘6�r�Fb��r�S*H�н�/���q�|���L�1}����J����h	u?�snt(�o`��V���rB�x $P�_��v4�;���h��5���q�Ʋ��	�� �K�>�hv(��0��gW��^�,P&�(��t�PZʂ"/�k�U�A��.�
I��ރ�	���+�?��>8�O&�({���SL�u(��0��t}pʄBR �l�B}�Ueq���$ׄBR ����AL�;p�\?�lL���Lh $PHh���3���"L_ۄ9�%	UҦM��4{�J�LQL[`�'@+��� �7��@Hn�I6�|my��Q(mYݼ�FLׂ2i����=���P�����p����j�&�(dn�F7�)�4�O��c%&뺬B(wcZ��(��)M
�|�rL���tK�(ӤR qL_���Q��&�(b+�a6���A��j�    IEND�B`�PK
      RZ���  �  /   images/7260fbed-8271-43c5-b1e8-f8e9900a221b.png�PNG

   IHDR  �      ��֗   gAMA  ���a    cHRM  z&  ��  �   ��  u0  �`  :�  p��Q<   bKGD ���̿   tIME�6���_  �IDATx��ܱM�P E�g+�^ �3K�Q�53�`�`��HP�q�o���ra��FI�                                                                                       ��T&X�&g���gg,(�6?�^[S�_m�< y@����$H�< y@��A����$H�< y@������$H�< y@����$H$H�< y@����$H�< y@� y@����$H�< y@��Ƀ���$H�< y@����$�$H�< y@����$H�<H� y@����$H�< y@��Ƀ���$H�< y@����$�$H�< y@����$H�<H�< y@����$H�< y@��A����$H�< y@������$H�< y@����$H$H�< y@����$H�< y��	@����$H�< y@������$H�< y@����$H$H�< y@����$H�< y�< y@����$H�< y@��Ƀ���$H�< y@����$�$H�< y@����$H�<H�< y@����$H�< y@� y����$H�< y@����$�$H�< y@����$H�<H�< y@����$H�< y@� y@����$H�< y@������$H�< y@����$H$H�< y@����$H�< y�< y@����$H�< y@��A�& ��$H�< y@����$H$H�< y@����$H�< y�< y@����$H�< y@��A����$H�< y@��������k6���&�^�}gg����ߋ��[۴�Z�uϯ���a�˛ $H�< y@����$H�< y�< y@��i�>�.�i�pN2                                     ��*��s����%��Ȼ�'w��������H$H�< y@����$H�< y�< y@�䁉[�ԇ bv&                                       8����νzȋ�������=�`�	@����$H�< y@������$H�<0��[�0xC                                                                                                                                          ���+b��0   %tEXtdate:create 2023-04-18T17:15:54+00:00SMK�   %tEXtdate:modify 2023-04-18T17:15:54+00:00"�=    IEND�B`�PK
      RZ�wp�&
  &
  /   images/e3aa425b-adcd-4ef1-9309-97e806748a2c.png�PNG

   IHDR  �      ��֗   gAMA  ���a   	pHYs  �  ��+   %tEXtdate:create 2023-04-18T17:15:54+00:00SMK�   %tEXtdate:modify 2023-04-18T17:15:54+00:00"�=  	fIDATx���!�Va���1�l�tW�&l&�f�=�Y��`uF NW܁#8�~��2s��<�N}�KߝB$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)�/8�{����a�$_�~^t�a^;'yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yHYN����qr�݋y>���y��r9�WC�ݫa?+����C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C�r���-��.����`�<�!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)�L��<�i���l�6�8�n������f��5IR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR����? bw.g�����9���<pM���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�H~���p���u��$���y:���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E��8�w�q·H~����-$yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)�#=Ng    IEND�B`�PK 
      RZ�9��n  �n                   cirkitFile.jsonPK 
      RZ                        &o  jsons/PK 
      RZ��                 Jo  jsons/user_defined.jsonPK 
      RZ                        ��  images/PK 
      RZuA�V� V� /             ��  images/61f598ae-58c3-4b7b-a0c5-99e4be3565c0.pngPK 
      RZ蓎�ɣ  ɣ  /             IH images/b240e25a-70ca-477b-8a45-be7a3295a83b.pngPK 
      RZX�U&: &: /             _� images/9bab9bed-0662-4eeb-a3ad-16a556afeca0.pngPK 
      RZ�7.-c&  c&  /             �& images/0291db46-fb1c-4fc7-8f6c-e1e807286f19.pngPK 
      RZ	��} } /             �M images/bbfae99c-8036-4c5e-89fd-a87441410720.pngPK 
      RZd��   �   /             ��	 images/a262aa33-74c4-460b-b0ad-c746896f6744.pngPK 
      RZ+L$��� �� /             ��	 images/d8ab57a1-5a79-4c55-bee7-02b60939cb6a.pngPK 
      RZ���͗  �  /             ˬ images/cc0ca695-66e1-46bc-a2f3-28706ce884b5.pngPK 
      RZ���  �  /             �� images/7260fbed-8271-43c5-b1e8-f8e9900a221b.pngPK 
      RZ�wp�&
  &
  /             �� images/e3aa425b-adcd-4ef1-9309-97e806748a2c.pngPK      �  '�   